// This is the unpowered netlist.
module ram_controller (CEN_all,
    GWEN_0,
    GWEN_1,
    GWEN_2,
    GWEN_3,
    GWEN_4,
    GWEN_5,
    GWEN_6,
    GWEN_7,
    WEb_ram,
    ram_enabled,
    rst,
    wb_clk_i,
    A_all,
    D_all,
    Q0,
    Q1,
    Q2,
    Q3,
    Q4,
    Q5,
    Q6,
    Q7,
    WEN_all,
    bus_in,
    bus_out,
    requested_addr);
 output CEN_all;
 output GWEN_0;
 output GWEN_1;
 output GWEN_2;
 output GWEN_3;
 output GWEN_4;
 output GWEN_5;
 output GWEN_6;
 output GWEN_7;
 input WEb_ram;
 input ram_enabled;
 input rst;
 input wb_clk_i;
 output [8:0] A_all;
 output [7:0] D_all;
 input [7:0] Q0;
 input [7:0] Q1;
 input [7:0] Q2;
 input [7:0] Q3;
 input [7:0] Q4;
 input [7:0] Q5;
 input [7:0] Q6;
 input [7:0] Q7;
 output [7:0] WEN_all;
 input [7:0] bus_in;
 output [7:0] bus_out;
 input [15:0] requested_addr;

 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \requested_addr_latch[0] ;
 wire \requested_addr_latch[10] ;
 wire \requested_addr_latch[11] ;
 wire \requested_addr_latch[12] ;
 wire \requested_addr_latch[13] ;
 wire \requested_addr_latch[14] ;
 wire \requested_addr_latch[15] ;
 wire \requested_addr_latch[1] ;
 wire \requested_addr_latch[2] ;
 wire \requested_addr_latch[3] ;
 wire \requested_addr_latch[4] ;
 wire \requested_addr_latch[5] ;
 wire \requested_addr_latch[6] ;
 wire \requested_addr_latch[7] ;
 wire \requested_addr_latch[8] ;
 wire \requested_addr_latch[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A4 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__B2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__B2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__C1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__A4 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__116__A4 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__B2 (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__B2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__C1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__A4 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A4 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__B2 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__B2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__C1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__A4 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__A4 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__B2 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__B2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__C1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A4 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A3 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__B (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__A4 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A1 (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A2 (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__B2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(\requested_addr_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(\requested_addr_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__I (.I(\requested_addr_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__I (.I(\requested_addr_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__I (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A4 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A1 (.I(\requested_addr_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A2 (.I(\requested_addr_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A2 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__A2 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A4 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__B2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__C1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__A4 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A4 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__B2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__C1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A4 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A4 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__B2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__C1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__A4 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A4 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__B2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__C1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__A4 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__D (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__D (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__D (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__D (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__D (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__D (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__D (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__D (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__D (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__D (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__D (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__D (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(Q1[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(Q1[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(Q1[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(Q1[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(Q1[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(Q1[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(Q1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(Q2[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(Q2[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(Q2[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Q0[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(Q2[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(Q2[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(Q2[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(Q2[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(Q2[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(Q3[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(Q3[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(Q3[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(Q3[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(Q3[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Q0[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(Q3[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(Q3[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(Q3[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(Q4[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(Q4[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(Q4[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(Q4[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(Q4[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(Q4[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(Q4[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(Q0[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(Q4[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(Q5[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(Q5[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(Q5[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(Q5[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(Q5[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(Q5[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(Q5[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(Q5[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(Q6[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(Q0[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(Q6[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(Q6[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(Q6[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(Q6[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(Q6[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(Q6[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(Q6[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(Q7[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(Q7[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(Q7[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(Q0[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(Q7[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(Q7[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(Q7[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(Q7[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(Q7[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(WEb_ram));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(Q0[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(ram_enabled));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(requested_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(requested_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(requested_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(requested_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(requested_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(Q0[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(requested_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(requested_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(requested_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(requested_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(requested_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(requested_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(requested_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(requested_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(requested_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(requested_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(Q0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(requested_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(Q1[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _106_ (.I(_004_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _107_ (.I(_025_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _108_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net52),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _109_ (.A1(_068_),
    .A2(_070_),
    .A3(_072_),
    .A4(_075_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _110_ (.A1(_060_),
    .A2(_061_),
    .B1(_065_),
    .B2(_076_),
    .ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _111_ (.I(net5),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _112_ (.A1(net21),
    .A2(_062_),
    .B1(_063_),
    .B2(net45),
    .C1(net61),
    .C2(_064_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _113_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net13),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _114_ (.A1(_053_),
    .A2(net29),
    .A3(_069_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _115_ (.A1(_055_),
    .A2(net37),
    .B(_071_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _116_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net53),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _117_ (.A1(_079_),
    .A2(_080_),
    .A3(_081_),
    .A4(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _118_ (.A1(_077_),
    .A2(_061_),
    .B1(_078_),
    .B2(_083_),
    .ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _119_ (.I(net6),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _120_ (.A1(net22),
    .A2(_062_),
    .B1(_063_),
    .B2(net46),
    .C1(net62),
    .C2(_064_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _121_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net14),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _122_ (.A1(_053_),
    .A2(net30),
    .A3(_069_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _123_ (.A1(_055_),
    .A2(net38),
    .B(_071_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _124_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net54),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _125_ (.A1(_086_),
    .A2(_087_),
    .A3(_088_),
    .A4(_089_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _126_ (.A1(_084_),
    .A2(_061_),
    .B1(_085_),
    .B2(_090_),
    .ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _127_ (.I(net7),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _128_ (.A1(net23),
    .A2(_062_),
    .B1(_063_),
    .B2(net47),
    .C1(net63),
    .C2(_064_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _129_ (.A1(_066_),
    .A2(_067_),
    .A3(_015_),
    .A4(net15),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _130_ (.A1(_038_),
    .A2(net31),
    .A3(_069_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _131_ (.A1(_035_),
    .A2(net39),
    .B(_071_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _132_ (.A1(_073_),
    .A2(_074_),
    .A3(_008_),
    .A4(net55),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _133_ (.A1(_093_),
    .A2(_094_),
    .A3(_095_),
    .A4(_096_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _134_ (.A1(_091_),
    .A2(_061_),
    .B1(_092_),
    .B2(_097_),
    .ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _135_ (.I(net8),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _136_ (.A1(net24),
    .A2(_018_),
    .B1(_026_),
    .B2(net48),
    .C1(net64),
    .C2(_030_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _137_ (.A1(_011_),
    .A2(_006_),
    .A3(_015_),
    .A4(net16),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _138_ (.A1(_038_),
    .A2(net32),
    .A3(_020_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _139_ (.A1(_035_),
    .A2(net40),
    .B(_023_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _140_ (.A1(_004_),
    .A2(_025_),
    .A3(_008_),
    .A4(net56),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _141_ (.A1(_100_),
    .A2(_101_),
    .A3(_102_),
    .A4(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _142_ (.A1(_098_),
    .A2(_009_),
    .B1(_099_),
    .B2(_104_),
    .ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _143_ (.A1(\requested_addr_latch[14] ),
    .A2(\requested_addr_latch[12] ),
    .A3(\requested_addr_latch[13] ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _144_ (.A1(net74),
    .A2(_105_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _145_ (.A1(net65),
    .A2(\requested_addr_latch[15] ),
    .A3(_000_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _146_ (.I(_001_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _147_ (.I(\requested_addr_latch[1] ),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _148_ (.I(_003_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _149_ (.I(\requested_addr_latch[0] ),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _150_ (.I(_005_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _151_ (.I(\requested_addr_latch[2] ),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _152_ (.I(_007_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _153_ (.A1(_004_),
    .A2(_006_),
    .A3(_008_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _154_ (.I(_009_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _155_ (.A1(_002_),
    .A2(_010_),
    .ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _156_ (.I(_003_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _157_ (.I(_011_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _158_ (.I(_006_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _159_ (.I(\requested_addr_latch[2] ),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _160_ (.I(_014_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _161_ (.I(_015_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _162_ (.I(_001_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _163_ (.A1(_012_),
    .A2(_013_),
    .A3(_016_),
    .A4(_017_),
    .ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _164_ (.A1(_011_),
    .A2(_005_),
    .A3(_007_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _165_ (.I(_018_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _166_ (.A1(_002_),
    .A2(_019_),
    .ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _167_ (.A1(\requested_addr_latch[1] ),
    .A2(\requested_addr_latch[0] ),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _168_ (.I(_020_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _169_ (.A1(_016_),
    .A2(_017_),
    .A3(_021_),
    .ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _170_ (.I(_008_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _171_ (.A1(_003_),
    .A2(_005_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _172_ (.I(_023_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _173_ (.A1(_022_),
    .A2(_017_),
    .A3(_024_),
    .ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _174_ (.I(_005_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _175_ (.A1(_003_),
    .A2(_025_),
    .A3(_014_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _176_ (.I(_026_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _177_ (.A1(_002_),
    .A2(_027_),
    .ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _178_ (.I(_004_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _179_ (.I(_025_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _180_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(_017_),
    .ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _181_ (.A1(_007_),
    .A2(_020_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _182_ (.I(_030_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _183_ (.A1(_002_),
    .A2(_031_),
    .ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _184_ (.I(net1),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _185_ (.A1(net17),
    .A2(_019_),
    .B1(_027_),
    .B2(net41),
    .C1(net57),
    .C2(_031_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _186_ (.I(_014_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _187_ (.I(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _188_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net9),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _189_ (.A1(_016_),
    .A2(net25),
    .A3(_021_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _190_ (.I(_034_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _191_ (.A1(_038_),
    .A2(net33),
    .B(_024_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _192_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net49),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _193_ (.A1(_036_),
    .A2(_037_),
    .A3(_039_),
    .A4(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _194_ (.A1(_032_),
    .A2(_010_),
    .B1(_033_),
    .B2(_041_),
    .ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _195_ (.I(net2),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _196_ (.A1(net18),
    .A2(_019_),
    .B1(_027_),
    .B2(net42),
    .C1(net58),
    .C2(_031_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _197_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net10),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _198_ (.A1(_016_),
    .A2(net26),
    .A3(_021_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _199_ (.A1(_038_),
    .A2(net34),
    .B(_024_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _200_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net50),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _201_ (.A1(_044_),
    .A2(_045_),
    .A3(_046_),
    .A4(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _202_ (.A1(_042_),
    .A2(_010_),
    .B1(_043_),
    .B2(_048_),
    .ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _203_ (.I(net3),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _204_ (.A1(net19),
    .A2(_019_),
    .B1(_027_),
    .B2(net43),
    .C1(net59),
    .C2(_031_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(_034_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _206_ (.A1(_012_),
    .A2(_013_),
    .A3(_051_),
    .A4(net11),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _207_ (.I(_015_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _208_ (.A1(_053_),
    .A2(net27),
    .A3(_021_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _209_ (.I(_034_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _210_ (.A1(_055_),
    .A2(net35),
    .B(_024_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _211_ (.I(_007_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _212_ (.A1(_028_),
    .A2(_029_),
    .A3(_057_),
    .A4(net51),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _213_ (.A1(_052_),
    .A2(_054_),
    .A3(_056_),
    .A4(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _214_ (.A1(_049_),
    .A2(_010_),
    .B1(_050_),
    .B2(_059_),
    .ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _215_ (.I(net4),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _216_ (.I(_009_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _217_ (.I(_018_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _218_ (.I(_026_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _219_ (.I(_030_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _220_ (.A1(net20),
    .A2(_062_),
    .B1(_063_),
    .B2(net44),
    .C1(net60),
    .C2(_064_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _221_ (.I(_011_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _222_ (.I(_006_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _223_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net12),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _224_ (.I(_020_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _225_ (.A1(_053_),
    .A2(net28),
    .A3(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _226_ (.I(_023_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _227_ (.A1(_055_),
    .A2(net36),
    .B(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _228_ (.D(net75),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _229_ (.D(net82),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _230_ (.D(net83),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _231_ (.D(net84),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _232_ (.D(net85),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _233_ (.D(net86),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _234_ (.D(net87),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _235_ (.D(net88),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _236_ (.D(net89),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _237_ (.D(net90),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _238_ (.D(net76),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _239_ (.D(net77),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _240_ (.D(net78),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _241_ (.D(net79),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _242_ (.D(net80),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _243_ (.D(net81),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _252_ (.I(net84),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _253_ (.I(net85),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _254_ (.I(net86),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _255_ (.I(net87),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _256_ (.I(net88),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _257_ (.I(net89),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _258_ (.I(net90),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _259_ (.I(net76),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _260_ (.I(net77),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(net91),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _262_ (.I(net66),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(net67),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _264_ (.I(net68),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _265_ (.I(net69),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _266_ (.I(net70),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(net71),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _268_ (.I(net72),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(net73),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(Q0[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(Q1[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(Q1[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(Q1[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(Q1[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(Q1[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(Q1[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(Q1[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(Q2[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(Q2[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(Q2[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(Q0[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(Q2[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(Q2[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(Q2[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(Q2[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(Q2[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(Q3[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(Q3[1]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(Q3[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(Q3[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(Q3[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(Q0[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(Q3[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(Q3[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(Q3[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(Q4[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(Q4[1]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(Q4[2]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(Q4[3]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(Q4[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(Q4[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(Q4[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(Q0[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(Q4[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input41 (.I(Q5[0]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(Q5[1]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(Q5[2]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(Q5[3]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(Q5[4]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(Q5[5]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(Q5[6]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(Q5[7]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(Q6[0]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(Q0[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(Q6[1]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input51 (.I(Q6[2]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(Q6[3]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input53 (.I(Q6[4]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(Q6[5]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input55 (.I(Q6[6]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input56 (.I(Q6[7]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input57 (.I(Q7[0]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input58 (.I(Q7[1]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input59 (.I(Q7[2]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(Q0[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input60 (.I(Q7[3]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input61 (.I(Q7[4]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(Q7[5]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input63 (.I(Q7[6]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input64 (.I(Q7[7]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input65 (.I(WEb_ram),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input66 (.I(bus_in[0]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(bus_in[1]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input68 (.I(bus_in[2]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input69 (.I(bus_in[3]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(Q0[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input70 (.I(bus_in[4]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input71 (.I(bus_in[5]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input72 (.I(bus_in[6]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input73 (.I(bus_in[7]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input74 (.I(ram_enabled),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input75 (.I(requested_addr[0]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input76 (.I(requested_addr[10]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input77 (.I(requested_addr[11]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(requested_addr[12]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(requested_addr[13]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(Q0[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(requested_addr[14]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(requested_addr[15]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(requested_addr[1]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(requested_addr[2]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(requested_addr[3]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(requested_addr[4]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input86 (.I(requested_addr[5]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input87 (.I(requested_addr[6]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input88 (.I(requested_addr[7]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input89 (.I(requested_addr[8]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(Q1[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input90 (.I(requested_addr[9]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(rst),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(A_all[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(CEN_all));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(D_all[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(D_all[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(D_all[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(D_all[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(D_all[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(D_all[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(D_all[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(D_all[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(GWEN_0));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(GWEN_1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(GWEN_2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(GWEN_3));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(GWEN_4));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(GWEN_5));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(GWEN_6));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(GWEN_7));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(A_all[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(A_all[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(A_all[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(A_all[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(A_all[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(A_all[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(A_all[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(A_all[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_133 (.ZN(net133));
 assign WEN_all[0] = net126;
 assign WEN_all[1] = net127;
 assign WEN_all[2] = net128;
 assign WEN_all[3] = net129;
 assign WEN_all[4] = net130;
 assign WEN_all[5] = net131;
 assign WEN_all[6] = net132;
 assign WEN_all[7] = net133;
endmodule

