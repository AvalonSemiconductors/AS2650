// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la_data_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [63:0] la_data_out;

 wire net146;
 wire net151;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net147;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net148;
 wire net116;
 wire net117;
 wire net118;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net149;
 wire net150;
 wire net119;
 wire net124;
 wire net120;
 wire net121;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net122;
 wire net123;
 wire net157;
 wire net130;
 wire net158;
 wire net131;
 wire net159;
 wire net132;
 wire net160;
 wire net133;
 wire net161;
 wire net134;
 wire net162;
 wire net135;
 wire net163;
 wire net136;
 wire net164;
 wire net137;
 wire net138;
 wire net165;
 wire net139;
 wire net166;
 wire net140;
 wire net167;
 wire net141;
 wire net168;
 wire net142;
 wire net169;
 wire net143;
 wire net170;
 wire net144;
 wire net171;
 wire net145;
 wire net172;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.alu_op[0] ;
 wire \as2650.alu_op[1] ;
 wire \as2650.alu_op[2] ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[12] ;
 wire \as2650.cycle[13] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ivec[0] ;
 wire \as2650.ivec[1] ;
 wire \as2650.ivec[2] ;
 wire \as2650.ivec[3] ;
 wire \as2650.ivec[4] ;
 wire \as2650.ivec[5] ;
 wire \as2650.ivec[6] ;
 wire \as2650.ivec[7] ;
 wire \as2650.last_intr ;
 wire \as2650.prefixed ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__I (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__I (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05854__I (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__I (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__I (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A1 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__A2 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__A2 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__A1 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__A3 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__B1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__B2 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__I (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A1 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A2 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__I (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__S (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__A1 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__A2 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__S0 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__S1 (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__A1 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__A2 (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__B1 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__B2 (.I(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__C1 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__A2 (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__I (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I0 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I3 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__S0 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A1 (.I(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A2 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__B2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__A2 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__I (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__S (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__S0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__S1 (.I(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A2 (.I(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__B2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__A2 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A1 (.I(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A2 (.I(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__S0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__A2 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__B2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__A2 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__B (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A2 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__B1 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__B2 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__B1 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A1 (.I(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__B1 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A3 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A2 (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A3 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__A2 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A2 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__A2 (.I(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__B1 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__B2 (.I(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A1 (.I(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A2 (.I(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A4 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A1 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A1 (.I(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__S0 (.I(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A2 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__B2 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A2 (.I(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A1 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A2 (.I(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__I (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A1 (.I(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__I (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__I (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__B2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A2 (.I(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__B (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__A2 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__I0 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__I (.I(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A2 (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A2 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__B2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A2 (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__A2 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__A1 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A2 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A3 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A1 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A2 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__I (.I(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A1 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A2 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__I (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__I (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__I (.I(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A2 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__A1 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__A2 (.I(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A1 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A2 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__I (.I(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__A2 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__A2 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__I (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__A1 (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A1 (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A2 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A3 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A1 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A2 (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__A2 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A2 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A2 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__I (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__I (.I(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__A2 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__I (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A2 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__I (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A2 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A2 (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A2 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A3 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A2 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A1 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A2 (.I(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A2 (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A3 (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__B2 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__C (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__I (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__I (.I(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__B (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__I (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A1 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__I (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__I (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__I (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__I (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__I (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__I (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A1 (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__I (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__A2 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__B1 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__B2 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__I (.I(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__I (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A1 (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A3 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A1 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A1 (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A2 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__I (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A2 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A1 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__B (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__I (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A2 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__I (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__I (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A2 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__I (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A2 (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__A1 (.I(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A1 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A3 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__I (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__B1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__B2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A2 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A2 (.I(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__I (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A2 (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A3 (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A4 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A1 (.I(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A3 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__I (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A3 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A1 (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__B (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__C (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__I (.I(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__I (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A1 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A3 (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__B (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A1 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A2 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A3 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A2 (.I(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__I (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A1 (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A2 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__I (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__I (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__I (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__I (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A1 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A3 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__A2 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__C (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__B (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__I (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__I (.I(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A1 (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A3 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A4 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__A1 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__A2 (.I(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__I (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__I (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A2 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A3 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A4 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__I (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__I (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A3 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A1 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__I (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A3 (.I(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A1 (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__I (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__I (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__I (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__I (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__I (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__I (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__B2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__B2 (.I(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A1 (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A2 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__B1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__B2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A3 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__I (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__I (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__I (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A2 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__I (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__I (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__I (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A1 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__B (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__C (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__I (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__I (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__I (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A1 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__I (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A2 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A4 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A1 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__I (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A1 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A4 (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A1 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__I (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__I (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A3 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06408__I (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__I (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__I (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A3 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A1 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__I (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A1 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__B2 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A2 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A2 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A3 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__I (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A1 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A2 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A1 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__I (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A1 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A2 (.I(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A1 (.I(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__B2 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A2 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__B (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A2 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__B2 (.I(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A1 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__I (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A2 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A2 (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__I (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__B (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A1 (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A3 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A4 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__I (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A1 (.I(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A4 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__I (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A3 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A3 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A4 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A1 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A1 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A3 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A1 (.I(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A2 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A3 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__B1 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__B2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A3 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__I (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A2 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A3 (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__B (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__I (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__I (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__I (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__I (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__I (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A1 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A2 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A1 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A2 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A4 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__I (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A2 (.I(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A2 (.I(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A3 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A4 (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A2 (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A3 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A1 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A2 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A2 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A1 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A2 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A2 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A4 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A2 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A1 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A3 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__I (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A1 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__I (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A1 (.I(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I1 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A1 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A2 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__I (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A2 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__B2 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A1 (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A2 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A2 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A2 (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__B2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__I (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A1 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A2 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__A1 (.I(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__I (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A1 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__B (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A1 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__I (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__I (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A1 (.I(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A3 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A2 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__I (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__I (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__I (.I(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A2 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A3 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__I (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__I (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__I (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A2 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A3 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A2 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A2 (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__I (.I(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A1 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A1 (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__B2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__I (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A2 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__B (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__B2 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__C (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__I (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A3 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__I (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A1 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A3 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A2 (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__B (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__I (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__I (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__I (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__I (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A2 (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A2 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A4 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__B (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A1 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__I (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A3 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A4 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__I (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__I (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__B1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__B2 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__B2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A2 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__I (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__I (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__I (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__I (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A3 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__B2 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A2 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__B2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__I (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A2 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__I (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A2 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__B (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__C (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__C (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A1 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__B2 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A2 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A2 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__I (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__B2 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A1 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__A1 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A1 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A2 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__A3 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__B (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__C (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__I (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__I (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I (.I(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__I (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__B1 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__B2 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A1 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__S (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A1 (.I(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__B2 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A3 (.I(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A4 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A2 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A3 (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A4 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__I (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__I (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__I (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__I (.I(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__B1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__I (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A2 (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A2 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__B1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__I (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A3 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A2 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__A1 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__B2 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A2 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__C2 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__I (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A1 (.I(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__I (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A1 (.I(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__B (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A3 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__I (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__B (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__C (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A2 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A2 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A2 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A2 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__B1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__B2 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A2 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__I (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A1 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A1 (.I(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__I (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__C2 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A2 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A2 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A1 (.I(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A2 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__B (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__B2 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__I (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A1 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A3 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__I (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A1 (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A4 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A2 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__I (.I(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A2 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__B (.I(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__I (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A1 (.I(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__B1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A2 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A2 (.I(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__C (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A2 (.I(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__B (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__C (.I(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__I1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A2 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__A2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A2 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A2 (.I(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A2 (.I(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__B2 (.I(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A1 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A2 (.I(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A3 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A2 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A2 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__A2 (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A1 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A1 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__B (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__B2 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A1 (.I(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A2 (.I(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A3 (.I(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A2 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A1 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A2 (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A3 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__B2 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A1 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A3 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__A1 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__B (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__C (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A4 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A1 (.I(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A2 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A3 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__I (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A2 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__B (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__I (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__I (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__I (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__I (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__I (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__I (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__C (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__I (.I(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__I (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__I (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__B (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__I (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__I (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__I (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__I (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__I (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__I (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__I (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__I (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__I (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__I (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A2 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__I (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A3 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__I (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__B (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__C (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__I (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A3 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A3 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__I (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A3 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A2 (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__B (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__I (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__I (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__I (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__I (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__I (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__B2 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__B2 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__I (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__I (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__I (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__C1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__C2 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__I (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__I (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__B (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__B2 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__C2 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__I (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__I (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__I (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__B1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__B2 (.I(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A1 (.I(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__B2 (.I(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A1 (.I(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__I (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__I (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__B2 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A1 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__B1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__B2 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__C1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__I (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__I (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A2 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__B1 (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__I (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__B1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__B2 (.I(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__I (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A2 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__B1 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A3 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A2 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__I (.I(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__I (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__I (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__I (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__B1 (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__B1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__B2 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__I (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__B1 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__B2 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__C2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__I (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__I (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__I (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__B1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__B1 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__I (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A2 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__B1 (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__B2 (.I(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__I (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__I (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__I (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__I (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__B1 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__B1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__I (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__I (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__I (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__B1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__C2 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__I (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__B (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A2 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__I (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__I (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__B1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__B1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__I (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__B1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A2 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__I (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__B1 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B1 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B2 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A2 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__B1 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__C2 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__B (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__B1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A2 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__B1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__B1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__B2 (.I(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__I (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__I (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__B1 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__I (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__I (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__B1 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A1 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A2 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__B1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__B2 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__B1 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__C1 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__B (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__B1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__I (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__B1 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__B1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__B1 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__I (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__B1 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__B1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__B2 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__B1 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__B2 (.I(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__C2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__B (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__B1 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__C1 (.I(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A2 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__B (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__B1 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A2 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__B1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A2 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__I (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A3 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__B2 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__I (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A3 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A1 (.I(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__B2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__B2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A1 (.I(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__I (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__B2 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__I (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__B1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__B2 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__I (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A2 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__B1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__B2 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__I (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__B1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__B2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A1 (.I(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__I (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__C (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__C (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__C (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__I (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__I (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A3 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__I (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__I (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__I (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__B (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__I (.I(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A1 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__I (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A1 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A2 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__I (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__I (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A3 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__I (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A1 (.I(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A2 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A1 (.I(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A1 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A2 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A1 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__I (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A1 (.I(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__I (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A3 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__I (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__I (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A1 (.I(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A1 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A4 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__B (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__C (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__I (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__B2 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__I (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A4 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__B (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__I (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__I (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__I (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__I (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__C (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__C (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__C (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__I (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__C (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__I (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__C (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__C (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__C (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A3 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__I (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__I (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__I (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__I (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__I (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__I (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__B (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__I (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__I (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__I (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__I (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__I (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__I (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__C (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__C (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A1 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__C (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__C (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__A1 (.I(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__I (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__I (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A3 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A2 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__B (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__B (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__B (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A1 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__I (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A2 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A1 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A3 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__I (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__B (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A1 (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A2 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A3 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A2 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A1 (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A4 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A2 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A2 (.I(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A3 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A1 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A3 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A4 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A3 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A3 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A4 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A1 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__I (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__I (.I(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A3 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A2 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A3 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__B (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A3 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__I (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A4 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__I (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__I (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__I (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__B2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A3 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__I (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__B (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__C (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A3 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__I (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A1 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A3 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__C (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__I (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__B (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__I (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__B (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A1 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A2 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A3 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A1 (.I(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__I (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A2 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A2 (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__I (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__C (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__B (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__I (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__I (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A1 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__I (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__I (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__I (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__I (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__I (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A2 (.I(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__I (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__I (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__I (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__I (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__I (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__I (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A1 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__C (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__I (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__B (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__B (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__I (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__B (.I(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__I (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__I (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A2 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__B (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__I (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__B (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__I (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A1 (.I(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__B (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__I (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__I (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__I (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__I (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__B (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__B (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__B (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A3 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__I (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A3 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A1 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__I (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__I (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__B (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A3 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A2 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__I (.I(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A3 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A3 (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A3 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__B (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A2 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__B1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__B2 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__B2 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A3 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A2 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__I (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__I (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__I (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A3 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__I (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A4 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__B (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A4 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A1 (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A2 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A3 (.I(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A2 (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__I (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__I (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__B2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A1 (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A2 (.I(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__I (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__I (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__I (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__I (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__I (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__I (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A3 (.I(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A4 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__I (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__I (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A3 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__B (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I (.I(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A2 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A3 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A1 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A2 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I0 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__I1 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__S (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__B (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__I (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__I (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__B1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__B2 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__B2 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__C1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__B (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__B1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__B2 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A2 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__B1 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__B2 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__B1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__B2 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__B1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__B (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__B1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__C (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__I (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__B (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__B2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B2 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__I (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B2 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__B2 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__I (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__I (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__B2 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__B1 (.I(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__B2 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__I (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__I (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A2 (.I(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__B1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__B2 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__B2 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B2 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__C2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A2 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A1 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__B1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__B2 (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__B1 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__C1 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__C2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__B1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__B2 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__C1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__C2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B2 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__B1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__B2 (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__B1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__B2 (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A2 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B1 (.I(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B2 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__I (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A4 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__I (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__I (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__B (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__I (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A3 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__I (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__B (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__I (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__I (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__A2 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__I (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__I (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A3 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__I (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__I (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__I (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__I (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__I (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__B (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__I (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__B (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__I (.I(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A3 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__I (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A3 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A3 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A1 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__B (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A3 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__I (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A3 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__B (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__B1 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I (.I(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__B1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__I (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A2 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__B (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A1 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__B (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__B1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__I (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A3 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__B2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__I0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__S (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__I0 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__S (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__B1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__I (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A1 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A1 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__I (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__I (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A1 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__I (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__I (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__I (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__I (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__I (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__I (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__I (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__I (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__B (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__B (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__I (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__I (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__I (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A1 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__B1 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A1 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A2 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A1 (.I(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__B1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A1 (.I(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A2 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A3 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__I (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__I (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__B (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__I (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__I (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__I (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A1 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__I (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__B1 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__I (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__I (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__I (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__I (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__I (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__I (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__I (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__I (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__I (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__I (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A3 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__I0 (.I(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__I1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__I0 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__I1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__I1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__I0 (.I(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__I1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__I (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__I (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__I (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__B (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__I (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A2 (.I(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__I (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__I (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__B (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__C (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__I (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__I (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__I (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__C (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A2 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A3 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__I (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__I (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A2 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__A2 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A1 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A1 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A2 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__C (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__B (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A3 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__I0 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A3 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A3 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__B (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A3 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A4 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__I (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A3 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A2 (.I(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A3 (.I(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A1 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A3 (.I(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A4 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A3 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A3 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A3 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A2 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A1 (.I(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A3 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__I (.I(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__B (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__I (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__I (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A1 (.I(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__B (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__I (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__B (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__B2 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__B1 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__B2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__C (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__I (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A2 (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__B1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__B2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__C (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A2 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__B (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__B2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__I (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__I (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__I (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A2 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A3 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__B2 (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A2 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__B1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__B2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__C (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__B (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__I (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__I0 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__I1 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__S (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A2 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__I (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__I (.I(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__I (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__B1 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__I (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A1 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__I (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__B (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A2 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__I (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__C1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__C2 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__I (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__I (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__B (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A2 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__A1 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A2 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A2 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A2 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__B (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__B (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__B (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__B2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__C (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__B2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__B2 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A1 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A2 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__I (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A1 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A2 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__B (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A2 (.I(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A3 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__B (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A1 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__I (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__B2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A3 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__I (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__B1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__C (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A2 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__B (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A2 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A1 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A2 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__B2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__I (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__I (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A2 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__I (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__I (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A2 (.I(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A2 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A2 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__B (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__B (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__I (.I(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__I (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__A2 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A1 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__B2 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A2 (.I(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__I (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__I (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B2 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__C1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__C2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A1 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__I (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__C (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__B (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__B (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__C (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__B (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A2 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__B (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__C (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B1 (.I(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__C2 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__B2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__B1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__I (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A2 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A2 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__B2 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A2 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__B1 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__B2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A2 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__B1 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__C (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__I (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__I (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__C (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__C (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__B (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A2 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__B (.I(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__B (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A2 (.I(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__I (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__I (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__B2 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__B (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__B2 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__I (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__I (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__B2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__A1 (.I(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__B (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A1 (.I(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__I (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__B2 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A2 (.I(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__C (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A1 (.I(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B2 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__C (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__I (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__I (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__B (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__B (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A2 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__B (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__B2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__B2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A2 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A2 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__B (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__B2 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__I (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__B2 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__B2 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__B2 (.I(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__A2 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A1 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A2 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__C (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A2 (.I(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__B2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__C (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A1 (.I(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__A2 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__B (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A3 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__B2 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__I (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__B (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A1 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__B2 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A2 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__A1 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__B2 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__B (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__C (.I(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__B2 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__B (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__I (.I(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__B (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A3 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A2 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A4 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A1 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A3 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A4 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__I (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__I (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A2 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__B (.I(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__C (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__A3 (.I(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A1 (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A3 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A4 (.I(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A3 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__B2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A1 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A3 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B3 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A2 (.I(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A3 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A4 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__A1 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A3 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A2 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A3 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A1 (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A2 (.I(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A3 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__B (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A4 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__C (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__C (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__I (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__C (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__B (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__C (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__A1 (.I(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A3 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A3 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__A2 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__I (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A3 (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A3 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__B (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__I0 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__I1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A1 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__B (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A1 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__I (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A2 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__B (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A3 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A2 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__B (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__C (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A2 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A3 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__B (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__C (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A2 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__B (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__C (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__I (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__C (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__C (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__I (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A1 (.I(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A2 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__I (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A2 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__B (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__I (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A2 (.I(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__B (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I0 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__B (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I0 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A2 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A2 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A2 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__A1 (.I(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__A2 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__B (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__I (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A2 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__I1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__I0 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A2 (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A3 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A4 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__I (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__I (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__I (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__B (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__C (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__B1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__B2 (.I(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__I (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__B1 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__B2 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__B1 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__B1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__B2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__B1 (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__B2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__I (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A2 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__B (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__A4 (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A3 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A4 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A3 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__I (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__I (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A1 (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A2 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__B1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__B2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__B1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__C1 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A1 (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A1 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__B2 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__B1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__B2 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__B2 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__A1 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__B1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A1 (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__A1 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A2 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__I0 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__S (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__A2 (.I(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A1 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A1 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A2 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__C (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__C (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A1 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__I (.I(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A2 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__C (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A2 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__B (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A1 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__B1 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__B2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__I (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__B2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__C (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__C (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__A1 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__A2 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__B (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__C (.I(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A2 (.I(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__C (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__I (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A1 (.I(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__I (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__I (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A2 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A2 (.I(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__I (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__I (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__A1 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__C2 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__A2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__B (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__B2 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__B1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__B2 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A1 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A2 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__B2 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__B2 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__B (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A2 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__C (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__C (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__I (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__I (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__I (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__I (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__I (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A2 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A3 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A2 (.I(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__B (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__I (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A1 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A2 (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__I (.I(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__A2 (.I(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__A2 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__I (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__B2 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__B2 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B1 (.I(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__B2 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B1 (.I(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__B2 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__B2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__B1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__B2 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__B1 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__C (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__B1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__B2 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__B1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__B2 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__B1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__B2 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__B1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__B2 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__B1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__B2 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__B1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__B2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__B1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__B2 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__B1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__B2 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__I (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A2 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__C (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A2 (.I(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__C (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A2 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A2 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__C (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A2 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__C (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__A2 (.I(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__B2 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__C (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A1 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A2 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__A2 (.I(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__I (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A2 (.I(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__C (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A1 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A2 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__B (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__I (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__A1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__B (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__B1 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__C (.I(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A2 (.I(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__C (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__B1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__B2 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__B1 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__B1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__B2 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__C1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__B (.I(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__B1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__B2 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__B1 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__B2 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__B1 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__B2 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__B1 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__B2 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__B (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__B1 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__C (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__C (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A2 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__I (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A2 (.I(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A2 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__B (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__C (.I(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A1 (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__C (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A2 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A2 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__B1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__B2 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__C2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A1 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__C (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A1 (.I(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A2 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__I (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__I (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__B2 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__I (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__B2 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__B2 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A1 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__B2 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__B2 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__B1 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__C (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__A1 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__C (.I(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__I (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__C (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A1 (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__I (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A1 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A2 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A2 (.I(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__B (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__C (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__I (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__B (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A1 (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A2 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__B (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__B1 (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__B2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A2 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A1 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__B2 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__I (.I(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__B (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A1 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__C (.I(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__C (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__I (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A2 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__C (.I(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A2 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__C (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A1 (.I(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A2 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A2 (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A2 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__B (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__A3 (.I(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A1 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A2 (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__B (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__C (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__C (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A1 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__C (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A2 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A2 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__C (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A1 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A2 (.I(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A2 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__I (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A2 (.I(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__C (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__A1 (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__B2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A1 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A2 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__C (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__C (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__I (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__B2 (.I(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A2 (.I(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__I (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A3 (.I(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__B (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__B (.I(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A1 (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__B (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__B1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__B (.I(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A1 (.I(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__B (.I(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__I1 (.I(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__S (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__B2 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__C (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__A2 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__C (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__C (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A1 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__A2 (.I(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__I (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__B1 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__B1 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__C (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__C (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A2 (.I(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__I (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__C (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A1 (.I(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A3 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__B2 (.I(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__C (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__I (.I(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A2 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__B (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__B1 (.I(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__B2 (.I(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A2 (.I(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__C (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__C (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__A2 (.I(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A2 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A2 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__A2 (.I(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__B1 (.I(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__C (.I(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__I (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__C (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A1 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__C (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A1 (.I(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__C (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__C (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A2 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A1 (.I(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__C (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__C (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__A2 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__C (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A2 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__C (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__B2 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__C (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A1 (.I(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__C (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A2 (.I(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A2 (.I(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__B (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__C (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A2 (.I(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A2 (.I(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__A1 (.I(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__B (.I(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__C (.I(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__B2 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__C (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__I (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A2 (.I(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__C (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A2 (.I(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__S (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__B2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__C (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A1 (.I(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__C (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__B (.I(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__C (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__B2 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__C (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__C (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__I (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__I (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A2 (.I(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__B (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__I (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__I (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__I (.I(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__I (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__I (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A2 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__B (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A2 (.I(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__I (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A2 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A2 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__I (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__C1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__C2 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__B1 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__B2 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A2 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__I (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__I (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__B1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__B2 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__I (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__B2 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__C (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__I (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__B1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__I (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__I (.I(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__B2 (.I(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__C (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__B (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A1 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__B1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__B2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A1 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__A2 (.I(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A2 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A1 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A1 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__B (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A2 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__B2 (.I(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__C (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A4 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__A1 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A2 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A3 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A2 (.I(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A3 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A1 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__I (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__B1 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__I (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__I (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__I (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A2 (.I(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A1 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A2 (.I(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A1 (.I(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__C (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A1 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A2 (.I(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__B (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A2 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__C (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A2 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__B (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__B (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__I (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__I (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__B1 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__B1 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__B2 (.I(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__C (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__I (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__B1 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__B2 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__C1 (.I(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__C2 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A2 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__I (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__B1 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__B2 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__C1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__B1 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__B2 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__C1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__C (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__B (.I(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__I (.I(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__B (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__A1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__B (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A1 (.I(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__B1 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__I (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A2 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__B2 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__C1 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__C2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__B1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__B2 (.I(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__C1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__C2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A1 (.I(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__B1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__C2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__I (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A2 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__B1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__C1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__C2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A1 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__B (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__B (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A1 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__B1 (.I(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__B2 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__C (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A2 (.I(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__C (.I(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A1 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__B (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__B (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__C (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A1 (.I(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B1 (.I(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__A1 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__B (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A2 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__B2 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__C1 (.I(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__C2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__I (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__B1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__B2 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__B1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__B2 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__C (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__B1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__B2 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__C2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A2 (.I(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A2 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__B1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__B2 (.I(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__C1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__C2 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A1 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__B (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__B1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__B2 (.I(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__C (.I(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A2 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A2 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__B (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A2 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A2 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__B (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__B1 (.I(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A2 (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__B1 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__C1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__C2 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A2 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__B1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__B2 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__C2 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__B1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__B2 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__C1 (.I(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__C2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__B1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__B2 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A1 (.I(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__B1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__B2 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__C (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B (.I(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A1 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__B1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A2 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__B (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A2 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__B (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__C (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__B1 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__B2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__C (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__I (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__B (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A2 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__B1 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__B2 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__C (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A2 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A2 (.I(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__B1 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__B2 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__C1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A1 (.I(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__C2 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__B1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__B2 (.I(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__C2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__B1 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A2 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A2 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__B (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__B (.I(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A2 (.I(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__B (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__I (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__B2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__B1 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__B1 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__B1 (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__B2 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__C1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__C2 (.I(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A2 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A2 (.I(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__B1 (.I(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__B2 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__C2 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__B2 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__C2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A2 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__B1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__B2 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__C1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__C2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__A1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__B1 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__B2 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__I (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A1 (.I(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A2 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A2 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A2 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A2 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A2 (.I(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A2 (.I(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__C (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__B1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__B2 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__C1 (.I(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__C2 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__B1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__B2 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__A1 (.I(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__C (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__B1 (.I(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__B2 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A2 (.I(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B1 (.I(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__C (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__B2 (.I(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__C1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__C2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A1 (.I(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A2 (.I(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__B (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__B (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A2 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__B1 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__B2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__B (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__B (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A2 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A4 (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A1 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__A2 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__B (.I(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__C (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A1 (.I(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__B (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__C (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A1 (.I(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A3 (.I(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__I (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__A1 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A1 (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__B (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__B (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A1 (.I(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__I (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A2 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__C (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__I (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__B (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__I (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__B (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__B (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A2 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__B (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A2 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__B (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A2 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__B (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A3 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A1 (.I(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__I (.I(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__A1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__B (.I(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__A2 (.I(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A1 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A1 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__A1 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__I (.I(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A1 (.I(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__A1 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A2 (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__A1 (.I(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__A2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A1 (.I(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__B1 (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A1 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A2 (.I(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A2 (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A2 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A3 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A2 (.I(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__C (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11500__B (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A2 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A1 (.I(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A1 (.I(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__A1 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__I (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__A1 (.I(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A2 (.I(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__A1 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A2 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__I (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__A1 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__I (.I(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__A2 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__A1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A2 (.I(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__A1 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__A2 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__A1 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__A2 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A1 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A1 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A2 (.I(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__B (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__C (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__B (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__C (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A1 (.I(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__B1 (.I(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__B2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A3 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A1 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A3 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__A1 (.I(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A1 (.I(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__A2 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__A2 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__C (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__A2 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__A1 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__B (.I(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A2 (.I(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__I (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11584__I (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__A2 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__A1 (.I(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__B2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__A2 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__A2 (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__I (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A2 (.I(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A2 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11597__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A1 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A1 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__A2 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__A1 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A2 (.I(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__B (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A1 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__B2 (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__C (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A1 (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__B2 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__C (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A1 (.I(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A3 (.I(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__A1 (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A1 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__A1 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__A1 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__B2 (.I(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__C (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A1 (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__B2 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__C (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A2 (.I(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A1 (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__B (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A1 (.I(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__B (.I(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__A2 (.I(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__B1 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A2 (.I(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__A1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__B (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__A1 (.I(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__B (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__A2 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__A2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A2 (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A1 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__B2 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A2 (.I(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__B1 (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__A2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A2 (.I(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__A1 (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__B (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A1 (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A2 (.I(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__B (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__B (.I(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__A2 (.I(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11656__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A3 (.I(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A1 (.I(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A2 (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A3 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__B (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11661__A1 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__C (.I(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__A1 (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__B (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__A1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__B (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__A1 (.I(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__A2 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__B2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__C (.I(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__A2 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A1 (.I(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__A1 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__B (.I(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__I0 (.I(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A1 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__B (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__A2 (.I(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__B (.I(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__CLK (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__D (.I(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__CLK (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__D (.I(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__CLK (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__D (.I(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12015__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__D (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__D (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__D (.I(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__D (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__D (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12041__D (.I(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__D (.I(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12043__D (.I(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12093__D (.I(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_170_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_171_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_171_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_172_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_173_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_173_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_175_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_176_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_178_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_179_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_179_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_181_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_181_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_185_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_187_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_188_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_189_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_189_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_191_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_191_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_192_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Left_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Left_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Left_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Left_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Left_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Left_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Left_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Left_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Left_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Left_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Left_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Left_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Left_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_694 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05842_ (.I(net5),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05843_ (.I(_05696_),
    .Z(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05844_ (.I(_05697_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05845_ (.I(_05698_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05846_ (.I(_05699_),
    .Z(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05847_ (.I(\as2650.ins_reg[4] ),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05848_ (.I(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05849_ (.I(_05702_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05850_ (.I(_05703_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05851_ (.I(net53),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05852_ (.I(\as2650.ins_reg[0] ),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05853_ (.I(_05706_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05854_ (.I(_05707_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05855_ (.I(_05708_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05856_ (.A1(_05705_),
    .A2(_05709_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05857_ (.I(_05709_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05858_ (.A1(net53),
    .A2(_05711_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05859_ (.I(net54),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05860_ (.I(\as2650.ins_reg[1] ),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05861_ (.I(_05714_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05862_ (.A1(_05713_),
    .A2(_05715_),
    .ZN(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05863_ (.I(net54),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05864_ (.I(_05714_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05865_ (.A1(_05717_),
    .A2(_05718_),
    .ZN(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05866_ (.A1(_05710_),
    .A2(_05712_),
    .A3(_05716_),
    .A4(_05719_),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05867_ (.I(\as2650.alu_op[2] ),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05868_ (.I(\as2650.alu_op[1] ),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05869_ (.I(_05722_),
    .ZN(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05870_ (.A1(_05721_),
    .A2(_05723_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05871_ (.I(_05724_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05872_ (.A1(_05709_),
    .A2(_05714_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05873_ (.I(_05726_),
    .Z(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05874_ (.A1(_05727_),
    .A2(_05720_),
    .ZN(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05875_ (.I(_05701_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05876_ (.I(_05721_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05877_ (.A1(_05730_),
    .A2(_05722_),
    .ZN(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05878_ (.A1(_05729_),
    .A2(_05731_),
    .ZN(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _05879_ (.A1(_05704_),
    .A2(_05720_),
    .A3(_05725_),
    .B1(_05728_),
    .B2(_05732_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05880_ (.I(_05729_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05881_ (.I(_05722_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05882_ (.A1(_05734_),
    .A2(_05735_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05883_ (.I(\as2650.r0[7] ),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05884_ (.I(_05737_),
    .Z(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05885_ (.A1(_05706_),
    .A2(\as2650.ins_reg[1] ),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05886_ (.I(_05739_),
    .Z(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05887_ (.I(_05740_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05888_ (.I(net51),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05889_ (.I(_05742_),
    .Z(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05890_ (.I(_05743_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05891_ (.I(_05744_),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05892_ (.I(_05745_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05893_ (.I(_05746_),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05894_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_05747_),
    .Z(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05895_ (.A1(_05706_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05896_ (.I(_05749_),
    .Z(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05897_ (.I(_05750_),
    .Z(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05898_ (.A1(\as2650.ins_reg[0] ),
    .A2(\as2650.ins_reg[1] ),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05899_ (.I(_05752_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05900_ (.I(_05753_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05901_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_05708_),
    .S1(_05747_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05902_ (.A1(_05738_),
    .A2(_05741_),
    .B1(_05748_),
    .B2(_05751_),
    .C1(_05754_),
    .C2(_05755_),
    .ZN(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05903_ (.I(_05756_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05904_ (.I(\as2650.r0[5] ),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05905_ (.I(_05758_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05906_ (.I(_05759_),
    .Z(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05907_ (.A1(_05760_),
    .A2(_05741_),
    .ZN(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05908_ (.I(_05746_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05909_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_05762_),
    .Z(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05910_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123[0][5] ),
    .I2(\as2650.r123_2[1][5] ),
    .I3(\as2650.r123_2[0][5] ),
    .S0(_05708_),
    .S1(_05762_),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05911_ (.A1(_05751_),
    .A2(_05763_),
    .B1(_05764_),
    .B2(_05754_),
    .ZN(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05912_ (.A1(_05761_),
    .A2(_05765_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05913_ (.I(\as2650.r0[4] ),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05914_ (.I(_05767_),
    .Z(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05915_ (.I(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05916_ (.I(_05740_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05917_ (.A1(_05769_),
    .A2(_05770_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05918_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_05746_),
    .Z(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05919_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_05707_),
    .S1(_05746_),
    .Z(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05920_ (.I(_05753_),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05921_ (.A1(_05750_),
    .A2(_05772_),
    .B1(_05773_),
    .B2(_05774_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05922_ (.A1(_05771_),
    .A2(_05775_),
    .ZN(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05923_ (.I(_05776_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05924_ (.I(\as2650.r0[3] ),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05925_ (.I(_05778_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05926_ (.I(_05779_),
    .ZN(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05927_ (.A1(_05708_),
    .A2(_05714_),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05928_ (.I(_05749_),
    .Z(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05929_ (.I(_05745_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05930_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_05783_),
    .Z(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05931_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_05707_),
    .S1(_05783_),
    .Z(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05932_ (.A1(_05782_),
    .A2(_05784_),
    .B1(_05785_),
    .B2(_05754_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05933_ (.A1(_05780_),
    .A2(_05781_),
    .B(_05786_),
    .ZN(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05934_ (.I(\as2650.r0[2] ),
    .Z(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05935_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_05745_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05936_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_05706_),
    .S1(_05745_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05937_ (.A1(_05788_),
    .A2(_05740_),
    .B1(_05789_),
    .B2(_05750_),
    .C1(_05790_),
    .C2(_05753_),
    .ZN(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05938_ (.I(_05791_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05939_ (.I(\as2650.r0[1] ),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05940_ (.I(_05793_),
    .Z(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05941_ (.I(_05743_),
    .Z(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05942_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_05795_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05943_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_05744_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05944_ (.A1(_05794_),
    .A2(_05739_),
    .B1(_05796_),
    .B2(_05749_),
    .C1(_05797_),
    .C2(_05752_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05945_ (.I(_05798_),
    .Z(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05946_ (.I(_05799_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05947_ (.I(\as2650.alu_op[0] ),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05948_ (.A1(\as2650.alu_op[2] ),
    .A2(\as2650.alu_op[1] ),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05949_ (.A1(_05701_),
    .A2(_05802_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05950_ (.I(\as2650.r0[0] ),
    .Z(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05951_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_05795_),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05952_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_05795_),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05953_ (.A1(_05804_),
    .A2(_05739_),
    .B1(_05805_),
    .B2(_05749_),
    .C1(_05806_),
    .C2(_05752_),
    .ZN(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05954_ (.I(_05807_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _05955_ (.A1(_05801_),
    .A2(_05803_),
    .A3(_05808_),
    .Z(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05956_ (.A1(_05792_),
    .A2(_05800_),
    .A3(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05957_ (.A1(_05777_),
    .A2(_05787_),
    .A3(_05810_),
    .ZN(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05958_ (.A1(_05766_),
    .A2(_05811_),
    .ZN(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05959_ (.A1(_05761_),
    .A2(_05765_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05960_ (.I(_05813_),
    .Z(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05961_ (.A1(_05771_),
    .A2(_05775_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05962_ (.I(_05815_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05963_ (.I(_05778_),
    .Z(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05964_ (.A1(_05817_),
    .A2(_05740_),
    .B1(_05784_),
    .B2(_05750_),
    .C1(_05785_),
    .C2(_05753_),
    .ZN(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05965_ (.I(_05818_),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05966_ (.I(_05791_),
    .Z(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05967_ (.I(_05799_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05968_ (.I(_05807_),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05969_ (.A1(_05721_),
    .A2(_05722_),
    .ZN(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05970_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.alu_op[0] ),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05971_ (.A1(_05823_),
    .A2(_05824_),
    .ZN(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05972_ (.A1(_05820_),
    .A2(_05821_),
    .A3(_05822_),
    .A4(_05825_),
    .Z(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05973_ (.A1(_05819_),
    .A2(_05826_),
    .Z(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05974_ (.A1(_05816_),
    .A2(_05827_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05975_ (.A1(_05814_),
    .A2(_05828_),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05976_ (.I(\as2650.r0[6] ),
    .Z(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05977_ (.I(_05830_),
    .Z(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05978_ (.I(_05831_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05979_ (.A1(_05832_),
    .A2(_05770_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05980_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_05762_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05981_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_05707_),
    .S1(_05762_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05982_ (.A1(_05751_),
    .A2(_05834_),
    .B1(_05835_),
    .B2(_05754_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05983_ (.A1(_05833_),
    .A2(_05836_),
    .Z(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05984_ (.I(_05837_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05985_ (.I0(_05812_),
    .I1(_05829_),
    .S(_05838_),
    .Z(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05986_ (.A1(_05757_),
    .A2(_05839_),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05987_ (.A1(_05833_),
    .A2(_05836_),
    .ZN(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05988_ (.I(_05841_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05989_ (.A1(_05812_),
    .A2(_05829_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05990_ (.A1(_00420_),
    .A2(_00421_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05991_ (.I(_05766_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05992_ (.A1(_05811_),
    .A2(_05828_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05993_ (.A1(_00423_),
    .A2(_00424_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05994_ (.I(_05819_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05995_ (.A1(_05810_),
    .A2(_05826_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05996_ (.A1(_00426_),
    .A2(_00427_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05997_ (.I(_05777_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05998_ (.I(_05787_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05999_ (.A1(_00430_),
    .A2(_05810_),
    .B(_05827_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06000_ (.A1(_00429_),
    .A2(_00431_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06001_ (.I(_05788_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06002_ (.I(_00433_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06003_ (.I(_00434_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06004_ (.I(_05781_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06005_ (.A1(_05782_),
    .A2(_05789_),
    .B1(_05790_),
    .B2(_05774_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06006_ (.A1(_00435_),
    .A2(_00436_),
    .B(_00437_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06007_ (.I(_05822_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06008_ (.A1(_00439_),
    .A2(_05825_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06009_ (.I(_05799_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06010_ (.I0(_05809_),
    .I1(_00440_),
    .S(_00441_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06011_ (.A1(_00438_),
    .A2(_00442_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06012_ (.I(_05804_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06013_ (.I(_00444_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06014_ (.A1(_00445_),
    .A2(_05741_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06015_ (.A1(_05782_),
    .A2(_05805_),
    .B1(_05806_),
    .B2(_05774_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06016_ (.A1(_00446_),
    .A2(_00447_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06017_ (.A1(_05803_),
    .A2(_00448_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06018_ (.A1(_05809_),
    .A2(_00440_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06019_ (.A1(_00441_),
    .A2(_00450_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06020_ (.A1(_00432_),
    .A2(_00443_),
    .A3(_00449_),
    .A4(_00451_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06021_ (.A1(_00428_),
    .A2(_00452_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06022_ (.A1(_05840_),
    .A2(_00422_),
    .A3(_00425_),
    .A4(_00453_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06023_ (.A1(_05736_),
    .A2(_00454_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06024_ (.A1(_05733_),
    .A2(_00455_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06025_ (.I(_00456_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06026_ (.I(_00457_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06027_ (.I(_00458_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06028_ (.I(\as2650.ins_reg[3] ),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06029_ (.A1(_00460_),
    .A2(_05729_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06030_ (.I(_00461_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06031_ (.I(_00462_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06032_ (.I(_00463_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06033_ (.I(\as2650.prefixed ),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06034_ (.I(_00465_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06035_ (.I(_05741_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06036_ (.I(\as2650.ins_reg[2] ),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06037_ (.I(_00460_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06038_ (.A1(_00468_),
    .A2(_00469_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06039_ (.I(_05802_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06040_ (.A1(_05701_),
    .A2(_05801_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06041_ (.A1(_00471_),
    .A2(_00472_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06042_ (.A1(_00470_),
    .A2(_00473_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06043_ (.A1(_00467_),
    .A2(_00474_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06044_ (.A1(net72),
    .A2(\as2650.cycle[0] ),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06045_ (.A1(_00475_),
    .A2(_00476_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06046_ (.A1(_00466_),
    .A2(_00477_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06047_ (.I(_05751_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06048_ (.I(_05721_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06049_ (.A1(_00480_),
    .A2(_05735_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06050_ (.I(_00469_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06051_ (.A1(_00482_),
    .A2(_05703_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06052_ (.A1(_00479_),
    .A2(_00481_),
    .A3(_00483_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06053_ (.I(_00484_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06054_ (.A1(_00478_),
    .A2(_00485_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06055_ (.A1(_05700_),
    .A2(_00459_),
    .A3(_00464_),
    .A4(_00486_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06056_ (.I(_00436_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _06057_ (.I(\as2650.ins_reg[2] ),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06058_ (.A1(_00489_),
    .A2(_00460_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06059_ (.I(_05729_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06060_ (.I(_05801_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06061_ (.A1(_00492_),
    .A2(_00471_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06062_ (.A1(_00491_),
    .A2(_00493_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06063_ (.A1(_00490_),
    .A2(_00494_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06064_ (.A1(_00488_),
    .A2(_00495_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06065_ (.I(net72),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06066_ (.A1(_00497_),
    .A2(\as2650.cycle[0] ),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06067_ (.I(_00498_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06068_ (.I(_00499_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06069_ (.A1(_00496_),
    .A2(_00500_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06070_ (.I(_00460_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06071_ (.A1(\as2650.prefixed ),
    .A2(_00502_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06072_ (.I(_00503_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06073_ (.A1(_00501_),
    .A2(_00504_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06074_ (.I(_00505_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06075_ (.I(_00468_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06076_ (.A1(_00507_),
    .A2(_05824_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06077_ (.A1(_05730_),
    .A2(_00508_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06078_ (.I(_00509_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06079_ (.A1(_05697_),
    .A2(_00510_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06080_ (.I(_00511_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06081_ (.I(_05698_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06082_ (.A1(_00513_),
    .A2(_00463_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06083_ (.I(_00465_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06084_ (.A1(_00515_),
    .A2(_00499_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06085_ (.A1(_00514_),
    .A2(_00516_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06086_ (.A1(_05726_),
    .A2(_05725_),
    .A3(_00461_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06087_ (.A1(_00507_),
    .A2(_00518_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06088_ (.I(_00519_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06089_ (.I(_00520_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06090_ (.I(_00521_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06091_ (.I(_05801_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06092_ (.A1(_00468_),
    .A2(_05702_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06093_ (.A1(_00523_),
    .A2(_00524_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06094_ (.A1(_05730_),
    .A2(_00525_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06095_ (.A1(_00482_),
    .A2(_00491_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06096_ (.A1(_00465_),
    .A2(_00527_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06097_ (.I(_00528_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06098_ (.I(_00529_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06099_ (.A1(net5),
    .A2(_00498_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06100_ (.I(_00531_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06101_ (.A1(_00526_),
    .A2(_00530_),
    .A3(_00532_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06102_ (.A1(_00506_),
    .A2(_00512_),
    .B1(_00517_),
    .B2(_00522_),
    .C(_00533_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06103_ (.I(\as2650.cycle[6] ),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06104_ (.I(_00535_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06105_ (.I(_00536_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06106_ (.I(_00537_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06107_ (.I(_00538_),
    .Z(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06108_ (.I(_00539_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06109_ (.I(_00540_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06110_ (.A1(_00487_),
    .A2(_00534_),
    .B(_00541_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06111_ (.I(net6),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06112_ (.I(_00543_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06113_ (.A1(_00544_),
    .A2(\as2650.cycle[1] ),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06114_ (.I(_00545_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06115_ (.I(_00546_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06116_ (.I(_00547_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06117_ (.I(net3),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06118_ (.I(_00549_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06119_ (.I(_00550_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06120_ (.I(_00551_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06121_ (.I(_00552_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06122_ (.I(_00553_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06123_ (.A1(_05699_),
    .A2(_00554_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06124_ (.A1(_00543_),
    .A2(\as2650.cycle[10] ),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06125_ (.A1(_00543_),
    .A2(\as2650.cycle[3] ),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06126_ (.I(net6),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06127_ (.I(_00558_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06128_ (.A1(_00559_),
    .A2(\as2650.cycle[1] ),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06129_ (.A1(_00557_),
    .A2(_00560_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06130_ (.A1(_00556_),
    .A2(_00561_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06131_ (.I(\as2650.addr_buff[7] ),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06132_ (.I(_00563_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06133_ (.I(_00564_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06134_ (.A1(_05699_),
    .A2(_00565_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06135_ (.A1(_00548_),
    .A2(_00555_),
    .B1(_00562_),
    .B2(_00566_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06136_ (.I(_05704_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06137_ (.I(_00568_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06138_ (.I(_00569_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06139_ (.I(_00570_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06140_ (.I(\as2650.cycle[9] ),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06141_ (.A1(_00559_),
    .A2(\as2650.cycle[2] ),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06142_ (.I(_00573_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06143_ (.I(_00574_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06144_ (.I(_00544_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06145_ (.A1(_00576_),
    .A2(\as2650.cycle[10] ),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06146_ (.I(_00577_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06147_ (.I(_00578_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06148_ (.I(_00561_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06149_ (.A1(_05698_),
    .A2(_00579_),
    .A3(_00580_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06150_ (.A1(_00571_),
    .A2(_00572_),
    .A3(_00575_),
    .A4(_00581_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06151_ (.I(\as2650.prefixed ),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06152_ (.A1(_00583_),
    .A2(_05703_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06153_ (.A1(_00499_),
    .A2(_00584_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06154_ (.A1(_00558_),
    .A2(\as2650.cycle[13] ),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06155_ (.I(_00586_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06156_ (.I(\as2650.cycle[11] ),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06157_ (.A1(_00543_),
    .A2(_00588_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06158_ (.A1(_00587_),
    .A2(_00589_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06159_ (.I(_00590_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06160_ (.A1(_00475_),
    .A2(_00585_),
    .A3(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06161_ (.A1(_00567_),
    .A2(_00582_),
    .B(_00592_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06162_ (.I(_00475_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06163_ (.I(_00585_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06164_ (.I(_00587_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06165_ (.A1(_00594_),
    .A2(_00595_),
    .A3(_00596_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06166_ (.A1(_00558_),
    .A2(\as2650.cycle[11] ),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06167_ (.I(_00598_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06168_ (.A1(_00597_),
    .A2(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06169_ (.A1(_00600_),
    .A2(_00575_),
    .A3(_00581_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06170_ (.I(_00583_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06171_ (.A1(_00602_),
    .A2(_00476_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06172_ (.A1(_00461_),
    .A2(_00603_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06173_ (.I(_00604_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06174_ (.A1(_00594_),
    .A2(_00484_),
    .A3(_00596_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06175_ (.I(_00606_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06176_ (.A1(_00558_),
    .A2(\as2650.cycle[5] ),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06177_ (.I(_00608_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06178_ (.I(_00609_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06179_ (.A1(_00544_),
    .A2(\as2650.cycle[4] ),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06180_ (.I(_00611_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06181_ (.A1(_00605_),
    .A2(_00607_),
    .A3(_00610_),
    .A4(_00612_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06182_ (.A1(_00559_),
    .A2(\as2650.cycle[13] ),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06183_ (.I(_00614_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06184_ (.I(_00615_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06185_ (.A1(_05696_),
    .A2(_00599_),
    .A3(_00613_),
    .B1(_00533_),
    .B2(_00616_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06186_ (.I(_00524_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06187_ (.A1(_00480_),
    .A2(_05735_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06188_ (.A1(_00523_),
    .A2(_00619_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06189_ (.A1(_00618_),
    .A2(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06190_ (.A1(_00523_),
    .A2(_05823_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06191_ (.I(_00622_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06192_ (.A1(_00623_),
    .A2(_00618_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06193_ (.A1(_00621_),
    .A2(_00624_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06194_ (.I(_00625_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06195_ (.A1(_00510_),
    .A2(_00530_),
    .A3(_00532_),
    .A4(_00626_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06196_ (.I(_00596_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06197_ (.I(_05731_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06198_ (.A1(_00468_),
    .A2(_00491_),
    .A3(_00629_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06199_ (.I(_00630_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06200_ (.I(_00631_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06201_ (.A1(_00525_),
    .A2(_00628_),
    .A3(_00632_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06202_ (.I(_00489_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06203_ (.A1(_00634_),
    .A2(_05732_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06204_ (.I(_00635_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06205_ (.I(_00624_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06206_ (.A1(_00636_),
    .A2(_00637_),
    .B(_00530_),
    .C(_00532_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06207_ (.I(_00532_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06208_ (.I(_00466_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(_00634_),
    .A2(_00518_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06210_ (.I(_00641_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06211_ (.I(_00615_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06212_ (.A1(_00504_),
    .A2(_00621_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06213_ (.A1(_00640_),
    .A2(_00642_),
    .A3(_00643_),
    .B(_00644_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06214_ (.I(\as2650.cycle[0] ),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06215_ (.I(net7),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06216_ (.A1(_00647_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06217_ (.A1(_00646_),
    .A2(_00648_),
    .B(_00497_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06218_ (.A1(_05696_),
    .A2(_00649_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06219_ (.A1(_00639_),
    .A2(_00645_),
    .B(_00650_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06220_ (.A1(_00627_),
    .A2(_00633_),
    .B(_00638_),
    .C(_00651_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06221_ (.I(\as2650.cycle[5] ),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06222_ (.A1(_00544_),
    .A2(_00653_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06223_ (.I(_00654_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06224_ (.I(_00655_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06225_ (.A1(_00576_),
    .A2(\as2650.cycle[7] ),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06226_ (.A1(_00519_),
    .A2(_00615_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06227_ (.A1(_00576_),
    .A2(\as2650.cycle[12] ),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06228_ (.I(_00659_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06229_ (.A1(_00605_),
    .A2(_00658_),
    .A3(_00660_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06230_ (.A1(_05697_),
    .A2(_00656_),
    .A3(_00657_),
    .A4(_00661_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06231_ (.A1(_00617_),
    .A2(_00652_),
    .A3(_00662_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06232_ (.A1(_00601_),
    .A2(_00663_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06233_ (.I(\as2650.cycle[13] ),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06234_ (.I(net5),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06235_ (.I(_00537_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06236_ (.I(_00667_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(_00666_),
    .A2(_00668_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06238_ (.I(_00669_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06239_ (.I(_00507_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06240_ (.A1(_00671_),
    .A2(_00484_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06241_ (.I(_00672_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06242_ (.I(_00673_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06243_ (.I(_00674_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06244_ (.I(_00605_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06245_ (.I(_00584_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06246_ (.I(_00677_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06247_ (.I(_00492_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06248_ (.A1(_00679_),
    .A2(_00481_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06249_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06250_ (.I(_00681_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06251_ (.I(_00682_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06252_ (.I(_00683_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06253_ (.I(_00684_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06254_ (.A1(_05703_),
    .A2(_00680_),
    .A3(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06255_ (.A1(_00467_),
    .A2(_00686_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06256_ (.A1(_00528_),
    .A2(_00687_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06257_ (.I(_00476_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06258_ (.A1(_00689_),
    .A2(_00630_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06259_ (.A1(_00688_),
    .A2(_00690_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06260_ (.A1(_00618_),
    .A2(_00620_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06261_ (.A1(_00622_),
    .A2(_00618_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06262_ (.A1(_00692_),
    .A2(_00693_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06263_ (.A1(_00508_),
    .A2(_00694_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06264_ (.A1(_00691_),
    .A2(_00695_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06265_ (.I(_00470_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06266_ (.I(_00477_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06267_ (.A1(_00678_),
    .A2(_00696_),
    .B(_00697_),
    .C(_00698_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06268_ (.A1(_00675_),
    .A2(_00676_),
    .B(_00699_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06269_ (.A1(_00670_),
    .A2(_00700_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06270_ (.A1(_00493_),
    .A2(_00593_),
    .B1(_00664_),
    .B2(_00665_),
    .C(_00701_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(_00542_),
    .A2(_00702_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06272_ (.I(_00689_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06273_ (.I(_00703_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06274_ (.I(_00529_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06275_ (.I(_00608_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06276_ (.I(_00706_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06277_ (.I(_00707_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06278_ (.A1(_00704_),
    .A2(_00511_),
    .A3(_00705_),
    .A4(_00708_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06279_ (.A1(_00663_),
    .A2(_00709_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06280_ (.I(_00710_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06281_ (.A1(_00601_),
    .A2(_00711_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06282_ (.I(_00712_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06283_ (.A1(_00489_),
    .A2(_00484_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06284_ (.I(_00714_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06285_ (.A1(_00715_),
    .A2(_00628_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06286_ (.I(_00478_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06287_ (.I(_00642_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06288_ (.I(_00718_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06289_ (.I(_00719_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06290_ (.I(_00720_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06291_ (.A1(_00564_),
    .A2(_00654_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06292_ (.I(_00722_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06293_ (.A1(_00514_),
    .A2(_00717_),
    .A3(_00721_),
    .A4(_00723_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06294_ (.A1(_00716_),
    .A2(_00724_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06295_ (.A1(\as2650.cycle[12] ),
    .A2(_00713_),
    .B(_00725_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06296_ (.I(_00726_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06297_ (.A1(_00588_),
    .A2(_00712_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06298_ (.I(_00628_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06299_ (.I(_00728_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06300_ (.I(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06301_ (.I(\as2650.cycle[4] ),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06302_ (.I(_00731_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06303_ (.I(_00639_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06304_ (.A1(_00515_),
    .A2(_05734_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06305_ (.I(_00734_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06306_ (.I(_00735_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06307_ (.A1(_00732_),
    .A2(_00733_),
    .A3(_00736_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06308_ (.A1(_00495_),
    .A2(_00730_),
    .A3(_00737_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06309_ (.I(_00485_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06310_ (.I(_00739_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06311_ (.I(_00707_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06312_ (.I(_00741_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06313_ (.A1(_00517_),
    .A2(_00612_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06314_ (.A1(_00740_),
    .A2(_00730_),
    .A3(_00742_),
    .A4(_00743_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06315_ (.A1(_00727_),
    .A2(_00738_),
    .A3(_00744_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06316_ (.I(_05700_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06317_ (.I(\as2650.cycle[3] ),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06318_ (.A1(_00559_),
    .A2(_00746_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06319_ (.I(_00747_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06320_ (.A1(_00748_),
    .A2(_00560_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06321_ (.I(\as2650.cycle[10] ),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06322_ (.A1(_00750_),
    .A2(_00713_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06323_ (.A1(_00745_),
    .A2(_00592_),
    .A3(_00749_),
    .B(_00751_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06324_ (.A1(_00600_),
    .A2(_00581_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06325_ (.A1(_00572_),
    .A2(_00710_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06326_ (.A1(_00575_),
    .A2(_00752_),
    .B(_00753_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06327_ (.I(_05699_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06328_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06329_ (.I(_00648_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06330_ (.A1(_00497_),
    .A2(_00756_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06331_ (.I(_00576_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06332_ (.I(_00704_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06333_ (.I(_00759_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06334_ (.I(_00760_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06335_ (.A1(_00758_),
    .A2(_00761_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06336_ (.I(\as2650.cycle[8] ),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06337_ (.I(_00763_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06338_ (.I(_00764_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06339_ (.I(_00765_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06340_ (.I(_00766_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06341_ (.A1(_00646_),
    .A2(_00757_),
    .B1(_00762_),
    .B2(_00767_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06342_ (.A1(_00755_),
    .A2(_00768_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06343_ (.A1(_00610_),
    .A2(_00658_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06344_ (.A1(_00754_),
    .A2(_00660_),
    .A3(_00769_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06345_ (.A1(\as2650.cycle[7] ),
    .A2(_00713_),
    .B1(_00770_),
    .B2(_00676_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06346_ (.I(_00771_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06347_ (.I(\as2650.cycle[8] ),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06348_ (.I(_00772_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06349_ (.A1(_00666_),
    .A2(_00476_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06350_ (.A1(_00773_),
    .A2(_00774_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06351_ (.I(_00775_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06352_ (.A1(_00541_),
    .A2(_00650_),
    .B1(_00776_),
    .B2(_00758_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06353_ (.I(_00777_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06354_ (.I(_00653_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06355_ (.I(_00587_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06356_ (.A1(_00698_),
    .A2(_00672_),
    .A3(_00779_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06357_ (.I(_05734_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06358_ (.I(_00781_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06359_ (.I(_00782_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06360_ (.I(_00783_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06361_ (.I(_00784_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06362_ (.I(_00785_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06363_ (.I(_00671_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06364_ (.I(_00787_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06365_ (.I(_00502_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06366_ (.I(_00789_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06367_ (.I(_00790_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06368_ (.I(_00791_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06369_ (.A1(_00788_),
    .A2(_00792_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06370_ (.I(_05697_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06371_ (.I(_00794_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06372_ (.I(_00640_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06373_ (.I(_00796_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06374_ (.I(_00797_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06375_ (.I(_00798_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06376_ (.A1(_00786_),
    .A2(_00793_),
    .B(_00795_),
    .C(_00799_),
    .ZN(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06377_ (.I(_00684_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06378_ (.I(_00801_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06379_ (.I(_00802_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06380_ (.I(_05730_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06381_ (.I(_05735_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06382_ (.I(_00472_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06383_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06384_ (.I(_00807_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06385_ (.I(_00808_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06386_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06387_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06388_ (.A1(_00805_),
    .A2(_00467_),
    .A3(_00806_),
    .A4(_00811_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06389_ (.A1(_00804_),
    .A2(_00812_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06390_ (.A1(_00803_),
    .A2(_00813_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06391_ (.A1(_00594_),
    .A2(_00585_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06392_ (.I(_00815_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06393_ (.I(_00816_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06394_ (.A1(_00473_),
    .A2(_00803_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06395_ (.I(_00629_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06396_ (.A1(_00819_),
    .A2(_00806_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06397_ (.I(_00820_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06398_ (.A1(_00817_),
    .A2(_00669_),
    .A3(_00818_),
    .A4(_00821_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06399_ (.A1(_00780_),
    .A2(_00800_),
    .B1(_00814_),
    .B2(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06400_ (.I(_00482_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06401_ (.I(_00824_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06402_ (.I(_00825_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06403_ (.A1(_00826_),
    .A2(_00665_),
    .A3(_00717_),
    .A4(_00511_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06404_ (.A1(_00778_),
    .A2(_00711_),
    .B(_00823_),
    .C(_00827_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06405_ (.I(_00666_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06406_ (.I(_00828_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06407_ (.I(_00829_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06408_ (.I(_00549_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06409_ (.I(_00831_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06410_ (.I(_00832_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06411_ (.I(_00833_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06412_ (.I(_00834_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06413_ (.I(_00835_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06414_ (.I(_00603_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06415_ (.I(_00719_),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06416_ (.I(_00483_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06417_ (.I(_00839_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06418_ (.A1(_00507_),
    .A2(_00587_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06419_ (.I(_00841_),
    .Z(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06420_ (.A1(_00840_),
    .A2(_00842_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06421_ (.A1(_00717_),
    .A2(_00720_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06422_ (.A1(_00837_),
    .A2(_00838_),
    .A3(_00730_),
    .B1(_00843_),
    .B2(_00844_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06423_ (.A1(_00830_),
    .A2(_00836_),
    .A3(_00845_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06424_ (.I(_00715_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06425_ (.I(_00847_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06426_ (.I(_00848_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06427_ (.I(_00616_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06428_ (.A1(_00849_),
    .A2(_00850_),
    .A3(_00724_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06429_ (.A1(_00623_),
    .A2(_00593_),
    .B1(_00710_),
    .B2(_00732_),
    .C(_00851_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06430_ (.A1(_00846_),
    .A2(_00852_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(_00746_),
    .A2(_00712_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06432_ (.A1(_00817_),
    .A2(_00670_),
    .A3(_00793_),
    .B(_00853_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06433_ (.A1(\as2650.cycle[1] ),
    .A2(_00713_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06434_ (.A1(_00788_),
    .A2(_00826_),
    .A3(_00670_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06435_ (.A1(_00595_),
    .A2(_00855_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06436_ (.A1(_00854_),
    .A2(_00856_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06437_ (.I(_00795_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06438_ (.A1(_00565_),
    .A2(_00562_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06439_ (.A1(_00836_),
    .A2(_00548_),
    .B(_00858_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06440_ (.A1(\as2650.cycle[2] ),
    .A2(_00712_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06441_ (.A1(_00857_),
    .A2(_00592_),
    .A3(_00859_),
    .B(_00860_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06442_ (.A1(_00721_),
    .A2(_00676_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06443_ (.A1(\as2650.cycle[13] ),
    .A2(_00609_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06444_ (.I(_00862_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06445_ (.I(_00863_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06446_ (.A1(_00849_),
    .A2(_00670_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06447_ (.A1(_00566_),
    .A2(_00864_),
    .B1(_00865_),
    .B2(_00459_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06448_ (.I(_00550_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06449_ (.I(_00867_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06450_ (.I(_00868_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06451_ (.I(_00869_),
    .Z(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06452_ (.A1(_00828_),
    .A2(_00870_),
    .A3(_00845_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06453_ (.A1(_00597_),
    .A2(_00613_),
    .B(_00589_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06454_ (.I(_00496_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06455_ (.I(_00653_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06456_ (.I(_00874_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06457_ (.A1(_00875_),
    .A2(_00595_),
    .B1(_00737_),
    .B2(_00474_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06458_ (.A1(_00873_),
    .A2(_00850_),
    .A3(_00876_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06459_ (.I(_00636_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06460_ (.I(_00878_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06461_ (.I(_00655_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06462_ (.I(_00880_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06463_ (.A1(_00513_),
    .A2(_00881_),
    .A3(_00661_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06464_ (.I(_00594_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06465_ (.A1(_00883_),
    .A2(_00643_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06466_ (.I(_00480_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06467_ (.I(_00508_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06468_ (.A1(_00885_),
    .A2(_00886_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06469_ (.A1(_00887_),
    .A2(_00631_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06470_ (.A1(_00627_),
    .A2(_00884_),
    .A3(_00888_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06471_ (.I(_00535_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06472_ (.I(_00890_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06473_ (.I(_00891_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06474_ (.A1(_00568_),
    .A2(_00892_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06475_ (.A1(_00837_),
    .A2(_00893_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06476_ (.I(_00488_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06477_ (.I(_00811_),
    .Z(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06478_ (.A1(_00494_),
    .A2(_00896_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06479_ (.A1(_00895_),
    .A2(_00897_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06480_ (.A1(_00894_),
    .A2(_00898_),
    .B(_05698_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06481_ (.A1(_00646_),
    .A2(_00650_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06482_ (.A1(_00759_),
    .A2(_00511_),
    .A3(_00705_),
    .A4(_00881_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06483_ (.I(_00797_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06484_ (.A1(_00646_),
    .A2(_00665_),
    .A3(_00588_),
    .A4(_00750_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06485_ (.A1(\as2650.cycle[1] ),
    .A2(_00746_),
    .A3(_00903_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06486_ (.I(\as2650.cycle[6] ),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06487_ (.I(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06488_ (.A1(_00778_),
    .A2(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06489_ (.A1(\as2650.cycle[4] ),
    .A2(_00907_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06490_ (.A1(\as2650.cycle[2] ),
    .A2(_00572_),
    .A3(\as2650.cycle[12] ),
    .A4(\as2650.cycle[7] ),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06491_ (.A1(_00904_),
    .A2(_00908_),
    .A3(_00909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06492_ (.A1(_00902_),
    .A2(_00873_),
    .B(_00639_),
    .C(_00910_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06493_ (.A1(_00899_),
    .A2(_00900_),
    .A3(_00901_),
    .A4(_00911_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06494_ (.A1(_00657_),
    .A2(_00882_),
    .B(_00889_),
    .C(_00912_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06495_ (.A1(_00533_),
    .A2(_00730_),
    .A3(_00879_),
    .B(_00913_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06496_ (.A1(_00871_),
    .A2(_00872_),
    .A3(_00877_),
    .A4(_00914_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06497_ (.A1(_00629_),
    .A2(_00806_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06498_ (.I(_00916_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06499_ (.A1(_00788_),
    .A2(_00795_),
    .A3(_00506_),
    .A4(_00917_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06500_ (.A1(_05718_),
    .A2(_00685_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06501_ (.I(_00523_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06502_ (.A1(_00920_),
    .A2(_05732_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06503_ (.A1(_00919_),
    .A2(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06504_ (.A1(_05711_),
    .A2(_00922_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06505_ (.I(_00923_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06506_ (.A1(_00691_),
    .A2(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06507_ (.I(_00687_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06508_ (.I(_05709_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06509_ (.I(_05715_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06510_ (.A1(_00927_),
    .A2(_00928_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06511_ (.A1(_00929_),
    .A2(_00896_),
    .A3(_00921_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06512_ (.I(_00930_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06513_ (.I(_00931_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06514_ (.A1(_00919_),
    .A2(_00921_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06515_ (.A1(_05711_),
    .A2(_00933_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06516_ (.I(_00934_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06517_ (.I(_00935_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06518_ (.I(_00929_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06519_ (.A1(_00937_),
    .A2(_00686_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06520_ (.A1(_00932_),
    .A2(_00936_),
    .A3(_00938_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06521_ (.A1(_00717_),
    .A2(_00926_),
    .A3(_00939_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06522_ (.I(_00504_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06523_ (.I(_00941_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06524_ (.A1(_00920_),
    .A2(_05724_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06525_ (.A1(_00491_),
    .A2(_00943_),
    .A3(_00811_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06526_ (.A1(_00488_),
    .A2(_00944_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06527_ (.A1(_00499_),
    .A2(_00945_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06528_ (.A1(_05704_),
    .A2(_00920_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06529_ (.A1(_00629_),
    .A2(_00947_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06530_ (.A1(_05727_),
    .A2(_00803_),
    .A3(_00948_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06531_ (.A1(_00942_),
    .A2(_00946_),
    .A3(_00949_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06532_ (.A1(_05727_),
    .A2(_00944_),
    .A3(_00696_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06533_ (.I(_00465_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06534_ (.I(_00952_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06535_ (.A1(_00953_),
    .A2(_00926_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06536_ (.A1(_00927_),
    .A2(_00928_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06537_ (.A1(_00955_),
    .A2(_00944_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06538_ (.I(_00956_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06539_ (.A1(_00733_),
    .A2(_00954_),
    .B1(_00957_),
    .B2(_00516_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06540_ (.A1(_00774_),
    .A2(_00644_),
    .B(_00638_),
    .C(_00958_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06541_ (.I(_00812_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06542_ (.A1(_00804_),
    .A2(_00817_),
    .A3(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06543_ (.I(_00467_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06544_ (.A1(_00733_),
    .A2(_00736_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06545_ (.A1(_00962_),
    .A2(_00897_),
    .A3(_00821_),
    .A4(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06546_ (.A1(_00951_),
    .A2(_00959_),
    .A3(_00961_),
    .A4(_00964_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06547_ (.A1(_00925_),
    .A2(_00940_),
    .A3(_00950_),
    .A4(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06548_ (.A1(_00918_),
    .A2(_00966_),
    .B(_00541_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06549_ (.A1(_00861_),
    .A2(_00866_),
    .B(_00915_),
    .C(_00967_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06550_ (.I(net95),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06551_ (.I(_05747_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06552_ (.A1(_00968_),
    .A2(_00962_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06553_ (.I(_00590_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06554_ (.A1(\as2650.cycle[8] ),
    .A2(_00774_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06555_ (.I(_00971_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06556_ (.A1(_00734_),
    .A2(_00972_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06557_ (.I(_00556_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06558_ (.A1(_00573_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06559_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06560_ (.A1(_00976_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06561_ (.I(_00977_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06562_ (.A1(_00975_),
    .A2(_00978_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06563_ (.A1(\as2650.cycle[9] ),
    .A2(_00979_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06564_ (.A1(_00747_),
    .A2(_00545_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06565_ (.A1(_00981_),
    .A2(_00908_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06566_ (.A1(_00970_),
    .A2(_00973_),
    .A3(_00980_),
    .A4(_00982_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06567_ (.A1(_00969_),
    .A2(_00983_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06568_ (.I(_00920_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06569_ (.I(_00985_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06570_ (.A1(_00986_),
    .A2(_00471_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06571_ (.A1(_05781_),
    .A2(_00977_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06572_ (.I(_00988_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06573_ (.A1(_00896_),
    .A2(_00989_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06574_ (.A1(_00874_),
    .A2(_00987_),
    .A3(_00990_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06575_ (.A1(_00905_),
    .A2(_00586_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06576_ (.I(_00992_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06577_ (.A1(_00968_),
    .A2(_00973_),
    .A3(_00991_),
    .A4(_00993_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06578_ (.I(_05747_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06579_ (.A1(_00995_),
    .A2(_00436_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06580_ (.I(_00996_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06581_ (.A1(\as2650.cycle[6] ),
    .A2(_00586_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06582_ (.A1(_00503_),
    .A2(_00526_),
    .A3(_00971_),
    .A4(_00998_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06583_ (.A1(_00997_),
    .A2(_00999_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06584_ (.I(_01000_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06585_ (.A1(_00984_),
    .A2(_00994_),
    .A3(_01001_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06586_ (.A1(\as2650.cycle[8] ),
    .A2(_00905_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06587_ (.I(_01003_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06588_ (.A1(_00602_),
    .A2(_00531_),
    .A3(_01004_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06589_ (.A1(_00897_),
    .A2(_01005_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06590_ (.A1(_00969_),
    .A2(_01006_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06591_ (.I(_01007_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06592_ (.A1(_00531_),
    .A2(_01003_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06593_ (.A1(_01009_),
    .A2(_00996_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06594_ (.A1(_00602_),
    .A2(_00502_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06595_ (.A1(_00941_),
    .A2(_00694_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06596_ (.A1(_05736_),
    .A2(_01011_),
    .B(_01012_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06597_ (.A1(_01010_),
    .A2(_01013_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06598_ (.I(_00969_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06599_ (.A1(_00772_),
    .A2(_00531_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06600_ (.A1(_00584_),
    .A2(_01016_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06601_ (.I(_00588_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06602_ (.A1(_00653_),
    .A2(\as2650.cycle[4] ),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06603_ (.I(_01019_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06604_ (.A1(_00535_),
    .A2(_00614_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06605_ (.A1(_01018_),
    .A2(_00562_),
    .A3(_01020_),
    .A4(_01021_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06606_ (.I(\as2650.addr_buff[6] ),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06607_ (.I(\as2650.addr_buff[5] ),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06608_ (.A1(_01023_),
    .A2(_01024_),
    .ZN(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06609_ (.A1(_00563_),
    .A2(_01025_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06610_ (.A1(_01017_),
    .A2(_01022_),
    .A3(_01026_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06611_ (.A1(_01015_),
    .A2(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06612_ (.A1(_01002_),
    .A2(_01008_),
    .A3(_01014_),
    .A4(_01028_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06613_ (.A1(_00937_),
    .A2(_01029_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06614_ (.I(_01030_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06615_ (.I(_00994_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06616_ (.I(_00680_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06617_ (.I(_01033_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06618_ (.I(_05808_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06619_ (.I(_00681_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06620_ (.A1(\as2650.holding_reg[0] ),
    .A2(_00682_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06621_ (.A1(_01035_),
    .A2(_01036_),
    .B(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06622_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06623_ (.I(_01039_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06624_ (.A1(_05770_),
    .A2(_01039_),
    .B(_00444_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06625_ (.A1(_00447_),
    .A2(_01040_),
    .B(_01041_),
    .C(_00682_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06626_ (.I(\as2650.holding_reg[0] ),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06627_ (.A1(_01043_),
    .A2(_00807_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06628_ (.A1(_01038_),
    .A2(_01042_),
    .A3(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06629_ (.I0(_01043_),
    .I1(_01035_),
    .S(_00808_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06630_ (.I(_01042_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06631_ (.I(_01044_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06632_ (.A1(_01047_),
    .A2(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06633_ (.A1(_01046_),
    .A2(_01049_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06634_ (.A1(_01045_),
    .A2(_01050_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06635_ (.A1(net50),
    .A2(net88),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06636_ (.A1(_01051_),
    .A2(_01052_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06637_ (.A1(_01034_),
    .A2(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06638_ (.I(_05725_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06639_ (.I(_00619_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06640_ (.A1(_00985_),
    .A2(_00819_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06641_ (.I(_01057_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06642_ (.A1(_01055_),
    .A2(_01056_),
    .A3(_01058_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06643_ (.I(_01059_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06644_ (.I(_00620_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06645_ (.I(_01061_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06646_ (.I(_01045_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06647_ (.A1(_00679_),
    .A2(_01056_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06648_ (.A1(_01062_),
    .A2(_01063_),
    .B1(_01050_),
    .B2(_01064_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06649_ (.A1(_01060_),
    .A2(_01065_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06650_ (.I(_01057_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06651_ (.I(net50),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06652_ (.I(net88),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06653_ (.A1(_01046_),
    .A2(_01047_),
    .A3(_01048_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06654_ (.A1(_01047_),
    .A2(_01048_),
    .B(_01046_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06655_ (.A1(_01068_),
    .A2(_01069_),
    .B(_01070_),
    .C(_01071_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06656_ (.A1(_01068_),
    .A2(_01069_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06657_ (.A1(_00679_),
    .A2(_01055_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06659_ (.A1(_01051_),
    .A2(_01073_),
    .B(_01075_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06660_ (.A1(_01067_),
    .A2(_01051_),
    .B1(_01072_),
    .B2(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06661_ (.I(_01059_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06662_ (.A1(_01054_),
    .A2(_01066_),
    .A3(_01077_),
    .B1(_01038_),
    .B2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(_01032_),
    .A2(net80),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06664_ (.A1(_01015_),
    .A2(_00983_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06665_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06666_ (.A1(_00976_),
    .A2(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06667_ (.I(_00976_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06668_ (.A1(_01084_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06669_ (.A1(_01083_),
    .A2(_01085_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06670_ (.I(_01086_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06671_ (.I(_01087_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06672_ (.A1(_00448_),
    .A2(_01088_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06673_ (.I(_01028_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06674_ (.I(_05808_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06675_ (.I(\as2650.addr_buff[5] ),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06676_ (.A1(_01023_),
    .A2(_01092_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06677_ (.I(_01023_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06678_ (.A1(_01094_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06679_ (.A1(_01093_),
    .A2(_01095_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06680_ (.A1(_01091_),
    .A2(_01096_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06681_ (.I(_01097_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06682_ (.I(_00445_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06683_ (.I(_01099_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06684_ (.A1(_01100_),
    .A2(_01008_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06685_ (.I(_01009_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06686_ (.I(_00997_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06687_ (.A1(_00504_),
    .A2(_00624_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06688_ (.A1(_01102_),
    .A2(_01103_),
    .A3(_01104_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06689_ (.I(_01105_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06690_ (.I(_01068_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06691_ (.I(_05756_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06692_ (.I(_01108_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06693_ (.A1(_01107_),
    .A2(_01109_),
    .B(_01052_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06694_ (.I(_00441_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06695_ (.A1(_00583_),
    .A2(_00482_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06696_ (.A1(_01112_),
    .A2(_00692_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06697_ (.A1(_01113_),
    .A2(_01010_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06698_ (.I(net8),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06699_ (.I(_01115_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06700_ (.I(_01116_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(_00614_),
    .A2(_00971_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06702_ (.A1(_00906_),
    .A2(_00503_),
    .A3(_00526_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06703_ (.A1(_00997_),
    .A2(_01118_),
    .A3(_01119_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06704_ (.I(_01120_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(_01113_),
    .A2(_01010_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06706_ (.A1(_00449_),
    .A2(_01120_),
    .B(_01122_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06707_ (.A1(_01117_),
    .A2(_01121_),
    .B(_01123_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06708_ (.A1(_01111_),
    .A2(_01114_),
    .B(_01105_),
    .C(_01124_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06709_ (.A1(_00466_),
    .A2(_01102_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06710_ (.A1(_00818_),
    .A2(_01126_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06711_ (.A1(_01103_),
    .A2(_01127_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06712_ (.I(_01128_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06713_ (.A1(_01106_),
    .A2(_01110_),
    .B(_01125_),
    .C(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06714_ (.I(_01028_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06715_ (.A1(_01101_),
    .A2(_01130_),
    .B(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06716_ (.A1(_01090_),
    .A2(_01098_),
    .B(_01132_),
    .C(_01081_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06717_ (.I(_00994_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06718_ (.A1(_01081_),
    .A2(_01089_),
    .B(_01133_),
    .C(_01134_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06719_ (.A1(_01080_),
    .A2(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06720_ (.I(_01099_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06721_ (.I(_01137_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06722_ (.I(_01138_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06723_ (.I(_00968_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06724_ (.I(_01140_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06725_ (.I(_01005_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06726_ (.A1(_01141_),
    .A2(_00926_),
    .A3(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06727_ (.I(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06728_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06729_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_05742_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06730_ (.I(_01146_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06731_ (.I(_01147_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06732_ (.I(_01148_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06733_ (.I(_01149_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06734_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06735_ (.A1(_01139_),
    .A2(_01145_),
    .A3(_01151_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06736_ (.A1(_00794_),
    .A2(_01143_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06737_ (.A1(_01153_),
    .A2(_01030_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06738_ (.I(_01154_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(\as2650.r123[1][0] ),
    .A2(_01155_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06740_ (.A1(_01031_),
    .A2(_01136_),
    .B(_01152_),
    .C(_01156_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06741_ (.I(_01030_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06742_ (.I(_00994_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06743_ (.A1(_05725_),
    .A2(_00619_),
    .A3(_01057_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06744_ (.I(_01159_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_05800_),
    .A2(_00808_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06746_ (.A1(\as2650.holding_reg[1] ),
    .A2(_00809_),
    .B(_01161_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06747_ (.I(\as2650.holding_reg[1] ),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06748_ (.A1(_05782_),
    .A2(_05796_),
    .B1(_05797_),
    .B2(_05774_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06749_ (.A1(_01164_),
    .A2(_01040_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06750_ (.I(_05794_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06751_ (.A1(_01166_),
    .A2(_00988_),
    .B(_00807_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06752_ (.A1(_01163_),
    .A2(_00808_),
    .B1(_01165_),
    .B2(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06753_ (.I(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06754_ (.A1(_01162_),
    .A2(_01169_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06755_ (.A1(_01070_),
    .A2(_01072_),
    .A3(_01170_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06756_ (.A1(_01070_),
    .A2(_01072_),
    .B(_01170_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06757_ (.A1(_01075_),
    .A2(_01171_),
    .A3(_01172_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06758_ (.A1(\as2650.holding_reg[1] ),
    .A2(_00682_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06759_ (.A1(_05821_),
    .A2(_01036_),
    .B(_01174_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06760_ (.A1(_01175_),
    .A2(_01168_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06761_ (.A1(_01047_),
    .A2(_01048_),
    .B(_01038_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06762_ (.A1(_01177_),
    .A2(_01052_),
    .B(_01045_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06763_ (.A1(_01176_),
    .A2(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06764_ (.A1(_01176_),
    .A2(_01178_),
    .B(_00943_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06765_ (.A1(_01179_),
    .A2(_01180_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06766_ (.A1(_01175_),
    .A2(_01169_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06767_ (.A1(_01175_),
    .A2(_01169_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06768_ (.I(_01159_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06769_ (.A1(_01061_),
    .A2(_01182_),
    .B1(_01183_),
    .B2(_01064_),
    .C(_01184_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06770_ (.A1(_01067_),
    .A2(_01170_),
    .B(_01185_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06771_ (.A1(_01181_),
    .A2(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06772_ (.A1(_01160_),
    .A2(_01162_),
    .B1(_01173_),
    .B2(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06773_ (.I(_01021_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06774_ (.I(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06775_ (.A1(_01020_),
    .A2(_01017_),
    .A3(_01026_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06776_ (.I(_00974_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06777_ (.A1(_00599_),
    .A2(_01192_),
    .A3(_00580_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06778_ (.A1(_01015_),
    .A2(_01190_),
    .A3(_01191_),
    .A4(_01193_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06779_ (.I(_01194_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06780_ (.A1(_05798_),
    .A2(_05807_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06781_ (.A1(\as2650.addr_buff[6] ),
    .A2(_01092_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06782_ (.A1(_05822_),
    .A2(_01093_),
    .B(_01197_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06783_ (.A1(_01196_),
    .A2(_01198_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06784_ (.I(_01199_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06785_ (.I(_01166_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06786_ (.I(_01201_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06787_ (.I(_05792_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06788_ (.I(_01203_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06789_ (.I(_01122_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06790_ (.I(_00503_),
    .Z(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06791_ (.A1(_01206_),
    .A2(_00637_),
    .A3(_01010_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06792_ (.I(net9),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06793_ (.I(_01208_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06794_ (.I(_01209_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06795_ (.I(_01210_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06796_ (.A1(_00997_),
    .A2(_01118_),
    .A3(_01119_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06797_ (.I(_01122_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_00451_),
    .A2(_01212_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06799_ (.A1(_01211_),
    .A2(_01212_),
    .B(_01213_),
    .C(_01214_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06800_ (.A1(_01204_),
    .A2(_01205_),
    .B(_01207_),
    .C(_01215_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06801_ (.I(_00439_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06802_ (.A1(_01217_),
    .A2(_01106_),
    .B(_01128_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06803_ (.A1(_01202_),
    .A2(_01129_),
    .B1(_01216_),
    .B2(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06804_ (.A1(_01194_),
    .A2(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06805_ (.A1(\as2650.cycle[9] ),
    .A2(_00589_),
    .A3(_00981_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06806_ (.A1(_01020_),
    .A2(_01017_),
    .A3(_00979_),
    .A4(_01189_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06807_ (.A1(_01103_),
    .A2(_01221_),
    .A3(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06808_ (.A1(_01195_),
    .A2(_01200_),
    .B(_01220_),
    .C(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06809_ (.I(_01083_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06810_ (.A1(_00976_),
    .A2(_01082_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06811_ (.A1(_01091_),
    .A2(_01225_),
    .B(_01226_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06812_ (.A1(_01196_),
    .A2(_01227_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06813_ (.I(_01228_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06814_ (.A1(_01081_),
    .A2(_01229_),
    .B(_01134_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06815_ (.A1(_01224_),
    .A2(_01230_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06816_ (.A1(_01158_),
    .A2(_01188_),
    .B(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06817_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_05743_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06818_ (.I(_01233_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06819_ (.I(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06820_ (.I(_01235_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06821_ (.I(_01236_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06822_ (.A1(_01201_),
    .A2(_00445_),
    .A3(_01150_),
    .A4(_01237_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06823_ (.I(_01202_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06824_ (.I(_01239_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06825_ (.A1(_01240_),
    .A2(_01151_),
    .B1(_01237_),
    .B2(_01137_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06826_ (.A1(_01238_),
    .A2(_01241_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06827_ (.I(_01242_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06828_ (.I(_01144_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06829_ (.A1(\as2650.r123[1][1] ),
    .A2(_01155_),
    .B1(_01243_),
    .B2(_01244_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06830_ (.A1(_01157_),
    .A2(_01232_),
    .B(_01245_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06831_ (.I(_00434_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06832_ (.I(_01246_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06833_ (.I(_01007_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06834_ (.I(_01111_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06835_ (.I(_01207_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06836_ (.I(net10),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06837_ (.I(_01251_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06838_ (.I(_01252_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06839_ (.A1(_01253_),
    .A2(_01000_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06840_ (.A1(_00443_),
    .A2(_01000_),
    .B(_01213_),
    .C(_01254_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06841_ (.A1(_00430_),
    .A2(_01205_),
    .B(_01207_),
    .C(_01255_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06842_ (.A1(_01249_),
    .A2(_01250_),
    .B(_01256_),
    .C(_01008_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06843_ (.A1(_01247_),
    .A2(_01248_),
    .B(_01131_),
    .C(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06844_ (.I(_01093_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06845_ (.A1(_05820_),
    .A2(_05821_),
    .A3(_05822_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06846_ (.A1(_00441_),
    .A2(_00439_),
    .B(_05792_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06847_ (.A1(_01260_),
    .A2(_01261_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _06848_ (.A1(_01259_),
    .A2(_01262_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06849_ (.A1(_05791_),
    .A2(_05799_),
    .A3(_05808_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06850_ (.A1(_05800_),
    .A2(_01091_),
    .B(_05792_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06851_ (.A1(_01259_),
    .A2(_01095_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06852_ (.I(_00438_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06853_ (.A1(_01264_),
    .A2(_01197_),
    .A3(_01265_),
    .B1(_01266_),
    .B2(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06854_ (.A1(_01263_),
    .A2(net81),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06855_ (.A1(_01194_),
    .A2(_01269_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06856_ (.I(_00984_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06857_ (.A1(_01258_),
    .A2(_01270_),
    .B(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06858_ (.A1(_01264_),
    .A2(_01226_),
    .A3(_01265_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06859_ (.A1(_01203_),
    .A2(_01087_),
    .B1(_01262_),
    .B2(_01225_),
    .C(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06860_ (.I(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06861_ (.A1(_01271_),
    .A2(_01275_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06862_ (.A1(\as2650.holding_reg[2] ),
    .A2(_00683_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06863_ (.A1(_01203_),
    .A2(_00801_),
    .B(_01277_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06864_ (.I(_00986_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06865_ (.A1(_01279_),
    .A2(_00481_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06866_ (.A1(_01162_),
    .A2(_01169_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06867_ (.I(_01036_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06868_ (.I(_01040_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06869_ (.A1(_05770_),
    .A2(_01040_),
    .B(_00434_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06870_ (.A1(_00437_),
    .A2(_01283_),
    .B(_01284_),
    .C(_01036_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06871_ (.A1(_00438_),
    .A2(_01282_),
    .B(_01285_),
    .C(\as2650.holding_reg[2] ),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06872_ (.A1(\as2650.holding_reg[2] ),
    .A2(_00683_),
    .B(_01285_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06873_ (.A1(_01203_),
    .A2(_01282_),
    .B(_01277_),
    .C(_01287_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06874_ (.A1(_01286_),
    .A2(_01288_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06875_ (.A1(_01172_),
    .A2(_01281_),
    .B(_01289_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06876_ (.A1(_01172_),
    .A2(_01289_),
    .A3(_01281_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06877_ (.A1(_01280_),
    .A2(_01290_),
    .A3(_01291_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06878_ (.I(_01289_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06879_ (.A1(_01182_),
    .A2(_01179_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06880_ (.A1(_01289_),
    .A2(_01294_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06881_ (.A1(_01279_),
    .A2(_01056_),
    .A3(_01286_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06882_ (.A1(_01064_),
    .A2(_01288_),
    .B(_01296_),
    .C(_01184_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06883_ (.A1(_01067_),
    .A2(_01293_),
    .B1(_01295_),
    .B2(_01034_),
    .C(_01297_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06884_ (.A1(_01060_),
    .A2(_01278_),
    .B1(_01292_),
    .B2(_01298_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06885_ (.A1(_01032_),
    .A2(_01299_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06886_ (.A1(_01158_),
    .A2(_01272_),
    .A3(_01276_),
    .B(_01300_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06887_ (.I(_01154_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06888_ (.A1(_01201_),
    .A2(_01236_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06889_ (.A1(_00434_),
    .A2(_01150_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06890_ (.I(\as2650.r0[2] ),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06891_ (.A1(_01305_),
    .A2(_01234_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06892_ (.A1(_01166_),
    .A2(_01149_),
    .A3(_01306_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06893_ (.A1(_01303_),
    .A2(_01304_),
    .B(_01307_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06894_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(_05742_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06895_ (.I(_01309_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06896_ (.I(_01310_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06897_ (.I(_01311_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06898_ (.I(_01312_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06899_ (.A1(_00445_),
    .A2(_01313_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06900_ (.A1(_01308_),
    .A2(_01314_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06901_ (.A1(_01238_),
    .A2(_01315_),
    .Z(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06902_ (.A1(\as2650.r123[1][2] ),
    .A2(_01302_),
    .B1(_01316_),
    .B2(_01244_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06903_ (.A1(_01157_),
    .A2(_01301_),
    .B(_01317_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06904_ (.I(_01134_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06905_ (.I(_00809_),
    .Z(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06906_ (.A1(_05819_),
    .A2(_00809_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06907_ (.A1(\as2650.holding_reg[3] ),
    .A2(_01319_),
    .B(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06908_ (.I(_01321_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06909_ (.I(_05779_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06910_ (.A1(_01323_),
    .A2(_00988_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06911_ (.A1(_05786_),
    .A2(_01283_),
    .B(_01324_),
    .C(_00683_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06912_ (.A1(\as2650.holding_reg[3] ),
    .A2(_01282_),
    .B(_01325_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06913_ (.I(_01326_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06914_ (.A1(_01321_),
    .A2(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06915_ (.I(_01328_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06916_ (.A1(_01293_),
    .A2(_01294_),
    .B(_01286_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06917_ (.A1(_01329_),
    .A2(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06918_ (.A1(_01278_),
    .A2(_01287_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06919_ (.A1(_01290_),
    .A2(_01332_),
    .B(_01328_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06920_ (.A1(_01290_),
    .A2(_01329_),
    .A3(_01332_),
    .Z(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06921_ (.A1(_01074_),
    .A2(_01333_),
    .A3(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06922_ (.A1(_01322_),
    .A2(_01326_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06923_ (.A1(_00985_),
    .A2(_00885_),
    .A3(_00805_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06924_ (.A1(_01058_),
    .A2(_01336_),
    .B(_01337_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06925_ (.A1(_01322_),
    .A2(_01326_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06926_ (.A1(_01061_),
    .A2(_01336_),
    .B1(_01338_),
    .B2(_01339_),
    .C(_01184_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06927_ (.A1(_01033_),
    .A2(_01331_),
    .B(_01335_),
    .C(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06928_ (.I(_01341_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06929_ (.A1(_01160_),
    .A2(_01322_),
    .B(_01342_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06930_ (.I(_01223_),
    .Z(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06931_ (.I(_01204_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06932_ (.I(_01213_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06933_ (.I(net11),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06934_ (.I(_01347_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06935_ (.I(_01348_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06936_ (.A1(_00428_),
    .A2(_01212_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06937_ (.A1(_01349_),
    .A2(_01212_),
    .B(_01205_),
    .C(_01350_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06938_ (.A1(_00429_),
    .A2(_01346_),
    .B(_01250_),
    .C(_01351_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06939_ (.A1(_01345_),
    .A2(_01250_),
    .B(_01352_),
    .C(_01248_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06940_ (.I(_05780_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06941_ (.A1(_01354_),
    .A2(_01129_),
    .B1(_01027_),
    .B2(_01015_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06942_ (.I(_01259_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06943_ (.A1(_05787_),
    .A2(_01260_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06944_ (.A1(_05818_),
    .A2(_01264_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06945_ (.I(_01095_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06946_ (.A1(_00430_),
    .A2(_01266_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06947_ (.A1(_01356_),
    .A2(_01357_),
    .B1(_01358_),
    .B2(_01359_),
    .C(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06948_ (.I(_01361_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06949_ (.A1(_01353_),
    .A2(_01355_),
    .B1(_01362_),
    .B2(_01195_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06950_ (.I(_01085_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06951_ (.A1(_01364_),
    .A2(_01358_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06952_ (.A1(_00426_),
    .A2(_01087_),
    .B1(_01357_),
    .B2(_01225_),
    .C(_01365_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06953_ (.I(_01366_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(_01223_),
    .A2(_01367_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06955_ (.A1(_01344_),
    .A2(_01363_),
    .B(_01368_),
    .C(_01134_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06956_ (.A1(_01318_),
    .A2(_01343_),
    .B(_01369_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06957_ (.A1(_01238_),
    .A2(_01315_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06958_ (.A1(_05788_),
    .A2(_01236_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06959_ (.I(\as2650.r0[3] ),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06960_ (.I(_01373_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06961_ (.A1(_01374_),
    .A2(_01148_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(_01372_),
    .A2(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06963_ (.A1(_01374_),
    .A2(_01149_),
    .A3(_01306_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06964_ (.A1(_01376_),
    .A2(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06965_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(net51),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06966_ (.I(_01379_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06967_ (.I(_01380_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06968_ (.A1(_05794_),
    .A2(_05804_),
    .A3(_01312_),
    .A4(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06969_ (.I(_01382_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06970_ (.A1(_05794_),
    .A2(_01312_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06971_ (.I(_01381_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(_00444_),
    .A2(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06973_ (.A1(_01384_),
    .A2(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(_01383_),
    .A2(_01387_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06975_ (.A1(_01378_),
    .A2(_01388_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06976_ (.A1(_01303_),
    .A2(_01304_),
    .B(_01307_),
    .C(_01314_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06977_ (.A1(_01307_),
    .A2(_01390_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06978_ (.A1(_01389_),
    .A2(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06979_ (.A1(_01371_),
    .A2(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06980_ (.I(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06981_ (.A1(\as2650.r123[1][3] ),
    .A2(_01302_),
    .B1(_01394_),
    .B2(_01145_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06982_ (.A1(_01157_),
    .A2(_01370_),
    .B(_01395_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06983_ (.A1(_05818_),
    .A2(_05820_),
    .A3(_05821_),
    .A4(_01035_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06984_ (.A1(_05815_),
    .A2(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06985_ (.A1(_01259_),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06986_ (.A1(_05819_),
    .A2(_05820_),
    .A3(_05800_),
    .A4(_01035_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06987_ (.A1(_05776_),
    .A2(_01399_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06988_ (.A1(_01359_),
    .A2(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06989_ (.A1(_05816_),
    .A2(_01096_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06990_ (.A1(_01398_),
    .A2(_01401_),
    .A3(_01402_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06991_ (.I(_00430_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06992_ (.I(_01105_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06993_ (.I(net12),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06994_ (.I(_01406_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06995_ (.I(_01407_),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06996_ (.I(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06997_ (.A1(_01409_),
    .A2(_01121_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06998_ (.A1(_00432_),
    .A2(_01001_),
    .B(_01346_),
    .C(_01410_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06999_ (.I(_00423_),
    .Z(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07000_ (.I(_01412_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07001_ (.A1(_01413_),
    .A2(_01114_),
    .B(_01405_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07002_ (.I(_01128_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07003_ (.A1(_01404_),
    .A2(_01405_),
    .B1(_01411_),
    .B2(_01414_),
    .C(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07004_ (.I(_05768_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07005_ (.I(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07006_ (.I(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07007_ (.A1(_01419_),
    .A2(_01248_),
    .B(_01090_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07008_ (.A1(_01416_),
    .A2(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07009_ (.A1(_01103_),
    .A2(_01221_),
    .A3(_01222_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07010_ (.A1(_01195_),
    .A2(_01403_),
    .B(_01421_),
    .C(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07011_ (.I(_05816_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07012_ (.I(_01225_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07013_ (.A1(_01364_),
    .A2(_01400_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07014_ (.A1(_01424_),
    .A2(_01087_),
    .B1(_01397_),
    .B2(_01425_),
    .C(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07015_ (.I(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07016_ (.A1(_01081_),
    .A2(_01428_),
    .B(_01318_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07017_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00802_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07018_ (.A1(_01424_),
    .A2(_00802_),
    .B(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07019_ (.A1(_01322_),
    .A2(_01327_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07020_ (.A1(_05816_),
    .A2(_01319_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07021_ (.A1(\as2650.holding_reg[4] ),
    .A2(_01319_),
    .B(_01433_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07022_ (.I(_01282_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07023_ (.I(_01283_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07024_ (.A1(_01418_),
    .A2(_00989_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07025_ (.A1(_05775_),
    .A2(_01436_),
    .B(_01437_),
    .C(_00684_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07026_ (.A1(\as2650.holding_reg[4] ),
    .A2(_01435_),
    .B(_01438_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07027_ (.A1(_01434_),
    .A2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07028_ (.I(_01440_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07029_ (.A1(_01434_),
    .A2(_01439_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07030_ (.I(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07031_ (.A1(_01441_),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07032_ (.A1(_01333_),
    .A2(_01432_),
    .B(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07033_ (.I(_01444_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07034_ (.A1(_01333_),
    .A2(_01446_),
    .A3(_01432_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07035_ (.A1(_01280_),
    .A2(_01445_),
    .A3(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07036_ (.A1(_01339_),
    .A2(_01330_),
    .B(_01336_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07037_ (.A1(_01446_),
    .A2(_01449_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07038_ (.A1(_00943_),
    .A2(_01450_),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07039_ (.A1(_01064_),
    .A2(_01440_),
    .B1(_01443_),
    .B2(_01062_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07040_ (.A1(_01279_),
    .A2(_00819_),
    .A3(_01446_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07041_ (.A1(_01060_),
    .A2(_01451_),
    .A3(_01452_),
    .A4(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07042_ (.A1(_01078_),
    .A2(_01431_),
    .B1(_01448_),
    .B2(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07043_ (.I(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _07044_ (.A1(_01423_),
    .A2(_01429_),
    .B1(_01456_),
    .B2(_01318_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07045_ (.I(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07046_ (.I(_00995_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07047_ (.I(_00945_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07048_ (.A1(_01459_),
    .A2(_01460_),
    .A3(_01126_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07049_ (.A1(_01371_),
    .A2(_01392_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07050_ (.A1(_01389_),
    .A2(_01391_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07051_ (.I(\as2650.r123[0][4] ),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07052_ (.A1(_05783_),
    .A2(\as2650.r123_2[0][4] ),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07053_ (.A1(_05783_),
    .A2(_01464_),
    .B(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07054_ (.I(_01466_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07055_ (.A1(_00444_),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07056_ (.A1(_01377_),
    .A2(_01468_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07057_ (.A1(_01376_),
    .A2(_01377_),
    .A3(_01382_),
    .A4(_01387_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07058_ (.A1(_05767_),
    .A2(_05778_),
    .A3(_01148_),
    .A4(_01235_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07059_ (.A1(_05769_),
    .A2(_01149_),
    .B1(_01236_),
    .B2(_05817_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07060_ (.A1(_01471_),
    .A2(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07061_ (.I(_01380_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07062_ (.A1(\as2650.r0[2] ),
    .A2(_05793_),
    .A3(_01310_),
    .A4(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07063_ (.I(_01475_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07064_ (.A1(_01383_),
    .A2(_01476_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07065_ (.A1(_00433_),
    .A2(_01313_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07066_ (.A1(\as2650.r0[1] ),
    .A2(_01474_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07067_ (.A1(_01383_),
    .A2(_01476_),
    .B1(_01478_),
    .B2(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07068_ (.A1(_01477_),
    .A2(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07069_ (.A1(_01470_),
    .A2(_01473_),
    .A3(_01481_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07070_ (.A1(_01469_),
    .A2(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07071_ (.A1(_01463_),
    .A2(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07072_ (.A1(_01462_),
    .A2(_01484_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07073_ (.A1(_01461_),
    .A2(_01485_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07074_ (.A1(\as2650.r123[1][4] ),
    .A2(_01155_),
    .B(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07075_ (.A1(_01157_),
    .A2(_01458_),
    .B(_01487_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07076_ (.A1(_05777_),
    .A2(_01396_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07077_ (.A1(_05814_),
    .A2(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07078_ (.A1(_05777_),
    .A2(_01399_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07079_ (.A1(_00423_),
    .A2(_01490_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07080_ (.A1(_01412_),
    .A2(_01088_),
    .B1(_01489_),
    .B2(_01425_),
    .C1(_01491_),
    .C2(_01364_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07081_ (.I(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07082_ (.A1(_01344_),
    .A2(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07083_ (.I(_05760_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07084_ (.I(_01495_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07085_ (.I(_01424_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07086_ (.I(net1),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07087_ (.I(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07088_ (.I(_01499_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07089_ (.I(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(_01501_),
    .A2(_01120_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07091_ (.A1(_00425_),
    .A2(_01000_),
    .B(_01213_),
    .C(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07092_ (.A1(_00420_),
    .A2(_01346_),
    .B(_01207_),
    .C(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07093_ (.A1(_01497_),
    .A2(_01250_),
    .B(_01504_),
    .C(_01008_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07094_ (.A1(_01496_),
    .A2(_01248_),
    .B(_01090_),
    .C(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07095_ (.A1(_05814_),
    .A2(_01266_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07096_ (.A1(_01356_),
    .A2(_01489_),
    .B1(_01491_),
    .B2(_01359_),
    .C(_01507_),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07097_ (.I(_01508_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07098_ (.A1(_01195_),
    .A2(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07099_ (.A1(_01506_),
    .A2(_01510_),
    .B(_01344_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07100_ (.A1(\as2650.holding_reg[5] ),
    .A2(_01435_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07101_ (.A1(_00423_),
    .A2(_00801_),
    .B(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07102_ (.I(_01513_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07103_ (.I(\as2650.holding_reg[5] ),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07104_ (.A1(_05765_),
    .A2(_01283_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07105_ (.A1(_01495_),
    .A2(_00989_),
    .B(_01516_),
    .C(_01319_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07106_ (.A1(_01515_),
    .A2(_00810_),
    .B(_01517_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07107_ (.A1(_01513_),
    .A2(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07108_ (.A1(_01514_),
    .A2(_01518_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07109_ (.A1(_01519_),
    .A2(_01520_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07110_ (.A1(_01442_),
    .A2(_01449_),
    .B(_01441_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07111_ (.A1(_01521_),
    .A2(_01522_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07112_ (.A1(_01431_),
    .A2(_01439_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07113_ (.A1(_01445_),
    .A2(_01524_),
    .B(_01521_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07114_ (.A1(_01445_),
    .A2(_01521_),
    .A3(_01524_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07115_ (.A1(_01075_),
    .A2(_01525_),
    .A3(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07116_ (.A1(_01514_),
    .A2(_01518_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07117_ (.I(_01337_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07118_ (.A1(_01067_),
    .A2(_01528_),
    .B(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07119_ (.I(_01519_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07120_ (.A1(_01062_),
    .A2(_01528_),
    .B1(_01530_),
    .B2(_01531_),
    .C(_01160_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07121_ (.A1(_01034_),
    .A2(_01523_),
    .B(_01527_),
    .C(_01532_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07122_ (.A1(_01078_),
    .A2(_01514_),
    .B(_01533_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07123_ (.A1(_01032_),
    .A2(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07124_ (.A1(_01158_),
    .A2(_01494_),
    .A3(_01511_),
    .B(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07125_ (.A1(_01377_),
    .A2(_01468_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07126_ (.A1(_01473_),
    .A2(_01477_),
    .A3(_01480_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07127_ (.A1(_01477_),
    .A2(_01480_),
    .B(_01473_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07128_ (.A1(_01470_),
    .A2(_01538_),
    .A3(_01539_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07129_ (.A1(_01469_),
    .A2(_01482_),
    .B(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07130_ (.I(\as2650.r123[0][5] ),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07131_ (.A1(_05744_),
    .A2(\as2650.r123_2[0][5] ),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07132_ (.A1(_05795_),
    .A2(_01542_),
    .B(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07133_ (.A1(_05804_),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07134_ (.A1(_01471_),
    .A2(_01545_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07135_ (.A1(_01166_),
    .A2(_01467_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07136_ (.A1(_01546_),
    .A2(_01547_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07137_ (.A1(_01383_),
    .A2(_01476_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07138_ (.A1(_01473_),
    .A2(_01480_),
    .B(_01549_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07139_ (.A1(_05759_),
    .A2(_05767_),
    .A3(_01147_),
    .A4(_01234_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07140_ (.A1(_05759_),
    .A2(_01148_),
    .B1(_01235_),
    .B2(_05768_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07141_ (.A1(_01551_),
    .A2(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07142_ (.A1(_01305_),
    .A2(_01381_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07143_ (.A1(_01374_),
    .A2(_01312_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07144_ (.A1(_01554_),
    .A2(_01555_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07145_ (.A1(_01373_),
    .A2(_01305_),
    .A3(_01311_),
    .A4(_01474_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07146_ (.A1(_01475_),
    .A2(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07147_ (.A1(_01553_),
    .A2(_01556_),
    .A3(_01558_),
    .Z(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07148_ (.A1(_01556_),
    .A2(_01558_),
    .B(_01553_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07149_ (.A1(_01559_),
    .A2(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07150_ (.A1(_01548_),
    .A2(_01550_),
    .A3(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07151_ (.A1(_01537_),
    .A2(_01541_),
    .A3(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_01463_),
    .A2(_01483_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07153_ (.A1(_01462_),
    .A2(_01484_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(_01564_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07155_ (.A1(_01563_),
    .A2(_01566_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07156_ (.I(_01567_),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07157_ (.A1(\as2650.r123[1][5] ),
    .A2(_01302_),
    .B1(_01568_),
    .B2(_01145_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07158_ (.A1(_01031_),
    .A2(_01536_),
    .B(_01569_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07159_ (.I(_05814_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07160_ (.I(net2),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07161_ (.I(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07162_ (.I(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07163_ (.I(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07164_ (.I(_01574_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07165_ (.I(_01575_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07166_ (.A1(_01576_),
    .A2(_01121_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07167_ (.A1(_00422_),
    .A2(_01001_),
    .B(_01205_),
    .C(_01577_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07168_ (.I(_01109_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07169_ (.A1(_01579_),
    .A2(_01114_),
    .B(_01106_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07170_ (.A1(_01570_),
    .A2(_01405_),
    .B1(_01578_),
    .B2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07171_ (.I(_05832_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07172_ (.I(_01582_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07173_ (.A1(_01583_),
    .A2(_01129_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07174_ (.A1(_01415_),
    .A2(_01581_),
    .B(_01584_),
    .C(_01131_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07175_ (.A1(_05813_),
    .A2(_05776_),
    .A3(_01396_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07176_ (.A1(_05841_),
    .A2(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07177_ (.A1(_05813_),
    .A2(_05776_),
    .A3(_01399_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07178_ (.A1(_05837_),
    .A2(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07179_ (.A1(_01356_),
    .A2(_01587_),
    .B1(_01589_),
    .B2(_01359_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07180_ (.A1(_00420_),
    .A2(_01266_),
    .B(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07181_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07182_ (.A1(_01194_),
    .A2(_01592_),
    .B(_01223_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07183_ (.A1(_01585_),
    .A2(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07184_ (.I(_05838_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07185_ (.A1(_01595_),
    .A2(_01088_),
    .B1(_01587_),
    .B2(_01425_),
    .C1(_01589_),
    .C2(_01364_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07186_ (.I(_01596_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07187_ (.A1(_01271_),
    .A2(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07188_ (.A1(_01318_),
    .A2(_01594_),
    .A3(_01598_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07189_ (.A1(_05841_),
    .A2(_00810_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07190_ (.A1(\as2650.holding_reg[6] ),
    .A2(_01435_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07191_ (.A1(_01600_),
    .A2(_01601_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07192_ (.I(_01514_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07193_ (.A1(_01603_),
    .A2(_01518_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07194_ (.A1(_01600_),
    .A2(_01601_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07195_ (.A1(_01582_),
    .A2(_00989_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07196_ (.A1(_05836_),
    .A2(_01436_),
    .B(_01606_),
    .C(_00684_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07197_ (.A1(\as2650.holding_reg[6] ),
    .A2(_00685_),
    .B(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07198_ (.A1(_01605_),
    .A2(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07199_ (.A1(_01605_),
    .A2(_01608_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07200_ (.I(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07201_ (.A1(_01609_),
    .A2(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07202_ (.I(_01612_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07203_ (.A1(_01525_),
    .A2(_01604_),
    .B(_01613_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07204_ (.A1(_01525_),
    .A2(_01613_),
    .A3(_01604_),
    .ZN(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07205_ (.A1(_01075_),
    .A2(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07206_ (.A1(_01528_),
    .A2(_01522_),
    .B(_01531_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07207_ (.A1(_01613_),
    .A2(_01617_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07208_ (.A1(_01058_),
    .A2(_01609_),
    .B(_01529_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07209_ (.A1(_01062_),
    .A2(_01609_),
    .B1(_01610_),
    .B2(_01619_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07210_ (.A1(_01614_),
    .A2(_01616_),
    .B1(_01618_),
    .B2(_01033_),
    .C(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07211_ (.A1(_01160_),
    .A2(_01602_),
    .B(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07212_ (.A1(_01158_),
    .A2(_01622_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07213_ (.A1(_01599_),
    .A2(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07214_ (.A1(_01564_),
    .A2(_01565_),
    .B(_01563_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07215_ (.A1(_01541_),
    .A2(_01562_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07216_ (.A1(_01541_),
    .A2(_01562_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07217_ (.A1(_01537_),
    .A2(_01626_),
    .B(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07218_ (.I(_01544_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07219_ (.I(_01629_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07220_ (.I(_01630_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07221_ (.A1(_01099_),
    .A2(_01471_),
    .A3(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07222_ (.I(_01466_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07223_ (.I(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07224_ (.A1(_01201_),
    .A2(_01634_),
    .A3(_01546_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(_01632_),
    .A2(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07226_ (.A1(_01559_),
    .A2(_01560_),
    .B(_01550_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07227_ (.A1(_01550_),
    .A2(_01559_),
    .A3(_01560_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07228_ (.A1(_01548_),
    .A2(_01637_),
    .B(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07229_ (.A1(_05793_),
    .A2(_01544_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07230_ (.A1(_01551_),
    .A2(_01640_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07231_ (.A1(_00433_),
    .A2(_01466_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07232_ (.A1(_01641_),
    .A2(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07233_ (.A1(_01476_),
    .A2(_01557_),
    .B(_01559_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07234_ (.I(\as2650.r123[0][6] ),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(_05743_),
    .A2(\as2650.r123_2[0][6] ),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07236_ (.A1(_05744_),
    .A2(_01645_),
    .B(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07237_ (.A1(\as2650.r0[0] ),
    .A2(_01647_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07238_ (.A1(_05830_),
    .A2(_05758_),
    .A3(_01147_),
    .A4(_01233_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07239_ (.A1(_05831_),
    .A2(_01147_),
    .B1(_01234_),
    .B2(_05759_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07240_ (.A1(_01649_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07241_ (.A1(_01648_),
    .A2(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07242_ (.I(_01311_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07243_ (.A1(_05767_),
    .A2(_01380_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07244_ (.A1(_05779_),
    .A2(_01653_),
    .A3(_01554_),
    .A4(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07245_ (.A1(\as2650.r0[3] ),
    .A2(_01474_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07246_ (.A1(_05768_),
    .A2(_01653_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07247_ (.A1(_01656_),
    .A2(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07248_ (.A1(_05788_),
    .A2(_01385_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07249_ (.A1(\as2650.r0[4] ),
    .A2(_01379_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07250_ (.A1(_05817_),
    .A2(_01653_),
    .A3(_01659_),
    .A4(_01660_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07251_ (.A1(_01655_),
    .A2(_01658_),
    .A3(_01661_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07252_ (.A1(_01652_),
    .A2(_01662_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07253_ (.A1(_01643_),
    .A2(_01644_),
    .A3(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07254_ (.A1(_01639_),
    .A2(_01664_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07255_ (.A1(_01636_),
    .A2(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _07256_ (.A1(_01625_),
    .A2(_01628_),
    .A3(_01666_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07257_ (.A1(_01461_),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07258_ (.A1(\as2650.r123[1][6] ),
    .A2(_01155_),
    .B(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07259_ (.A1(_01031_),
    .A2(_01624_),
    .B(_01669_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07260_ (.I(_00420_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07261_ (.A1(_00833_),
    .A2(_01121_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07262_ (.A1(_05840_),
    .A2(_01001_),
    .B(_01346_),
    .C(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07263_ (.A1(_01107_),
    .A2(_00448_),
    .B(_01073_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07264_ (.A1(_01114_),
    .A2(_01673_),
    .B(_01106_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07265_ (.A1(_01670_),
    .A2(_01405_),
    .B1(_01672_),
    .B2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07266_ (.I(_05738_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07267_ (.I(_01676_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07268_ (.I(_01677_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07269_ (.A1(_01678_),
    .A2(_01415_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07270_ (.A1(_01415_),
    .A2(_01675_),
    .B(_01679_),
    .C(_01090_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07271_ (.A1(_05838_),
    .A2(_01586_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07272_ (.A1(_01108_),
    .A2(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07273_ (.A1(_05838_),
    .A2(_01588_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07274_ (.A1(_05757_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07275_ (.A1(_01197_),
    .A2(_01684_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07276_ (.A1(_01108_),
    .A2(_01096_),
    .B1(_01682_),
    .B2(_01356_),
    .C(_01685_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07277_ (.I(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07278_ (.A1(_01131_),
    .A2(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07279_ (.A1(_01271_),
    .A2(_01688_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07280_ (.A1(_01226_),
    .A2(_01684_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07281_ (.A1(_01108_),
    .A2(_01088_),
    .B1(_01682_),
    .B2(_01425_),
    .C(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07282_ (.I(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07283_ (.A1(_01680_),
    .A2(_01689_),
    .B1(_01692_),
    .B2(_01344_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07284_ (.A1(\as2650.holding_reg[7] ),
    .A2(_01435_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07285_ (.A1(_05757_),
    .A2(_00801_),
    .B(_01694_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(_05757_),
    .A2(_00977_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07287_ (.A1(_01676_),
    .A2(_00977_),
    .B(_01696_),
    .C(_00685_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07288_ (.A1(\as2650.holding_reg[7] ),
    .A2(_00810_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07289_ (.I(_01695_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07290_ (.A1(_01697_),
    .A2(_01698_),
    .B(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07291_ (.I(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(_01697_),
    .A2(_01698_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07293_ (.A1(_01695_),
    .A2(_01702_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07294_ (.I(_01703_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07295_ (.A1(_01701_),
    .A2(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07296_ (.I(_01705_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07297_ (.A1(_01531_),
    .A2(_01522_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07298_ (.A1(_01528_),
    .A2(_01609_),
    .A3(_01707_),
    .B(_01610_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07299_ (.A1(_01706_),
    .A2(_01708_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07300_ (.A1(_01602_),
    .A2(_01608_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07301_ (.A1(_01614_),
    .A2(_01710_),
    .B(_01706_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07302_ (.A1(_01614_),
    .A2(_01706_),
    .A3(_01710_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07303_ (.A1(_01074_),
    .A2(_01711_),
    .A3(_01712_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07304_ (.A1(_01058_),
    .A2(_01700_),
    .B(_01529_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07305_ (.A1(_01061_),
    .A2(_01700_),
    .B1(_01704_),
    .B2(_01714_),
    .C(_01184_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07306_ (.A1(_01033_),
    .A2(_01709_),
    .B(_01713_),
    .C(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07307_ (.A1(_01060_),
    .A2(_01695_),
    .B(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07308_ (.I0(_01693_),
    .I1(_01717_),
    .S(_01032_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07309_ (.A1(_01628_),
    .A2(_01666_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07310_ (.A1(_01628_),
    .A2(_01666_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07311_ (.A1(_01625_),
    .A2(_01719_),
    .B(_01720_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07312_ (.I(_01636_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07313_ (.A1(_01549_),
    .A2(_01538_),
    .B(_01561_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07314_ (.A1(_01548_),
    .A2(_01723_),
    .A3(_01637_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(_01638_),
    .A2(_01724_),
    .B(_01664_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07316_ (.A1(_01722_),
    .A2(_01665_),
    .B(_01725_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07317_ (.I(_01640_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07318_ (.A1(_01641_),
    .A2(_01642_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07319_ (.A1(_01551_),
    .A2(_01727_),
    .B(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07320_ (.A1(_01644_),
    .A2(_01663_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07321_ (.A1(_01644_),
    .A2(_01663_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07322_ (.A1(_01643_),
    .A2(_01730_),
    .B(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07323_ (.A1(_01648_),
    .A2(_01649_),
    .A3(_01650_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07324_ (.A1(_01649_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07325_ (.A1(_00433_),
    .A2(_01629_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07326_ (.A1(_01734_),
    .A2(_01735_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07327_ (.A1(_05779_),
    .A2(_01633_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07328_ (.A1(_01736_),
    .A2(_01737_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07329_ (.A1(_01652_),
    .A2(_01655_),
    .A3(_01658_),
    .A4(_01661_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07330_ (.A1(_01661_),
    .A2(_01739_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07331_ (.A1(_05793_),
    .A2(_01647_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(_05830_),
    .A2(_01233_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07333_ (.A1(\as2650.r0[7] ),
    .A2(_01146_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07334_ (.A1(_01742_),
    .A2(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07335_ (.A1(_01741_),
    .A2(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07336_ (.A1(_01373_),
    .A2(_01311_),
    .A3(_01654_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07337_ (.A1(_05758_),
    .A2(_01309_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07338_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_05742_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07339_ (.A1(\as2650.r0[0] ),
    .A2(_01748_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07340_ (.A1(_01660_),
    .A2(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07341_ (.A1(_01747_),
    .A2(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07342_ (.A1(_01746_),
    .A2(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07343_ (.A1(_01745_),
    .A2(_01752_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07344_ (.A1(_01740_),
    .A2(_01753_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07345_ (.A1(_01732_),
    .A2(_01738_),
    .A3(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07346_ (.A1(_01729_),
    .A2(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07347_ (.A1(_01721_),
    .A2(_01726_),
    .A3(_01756_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07348_ (.I(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07349_ (.A1(\as2650.r123[1][7] ),
    .A2(_01302_),
    .B1(_01758_),
    .B2(_01145_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07350_ (.A1(_01031_),
    .A2(_01718_),
    .B(_01759_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07351_ (.I(_01069_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07352_ (.I(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07353_ (.A1(_00488_),
    .A2(_00802_),
    .A3(_00916_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07354_ (.A1(_00515_),
    .A2(_00971_),
    .A3(_01762_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07355_ (.I(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07356_ (.I(_01764_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07357_ (.I(net59),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07358_ (.I(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07359_ (.I(net89),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07360_ (.A1(_01767_),
    .A2(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07361_ (.I(_01769_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07362_ (.I(net70),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07363_ (.I(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07364_ (.A1(_01772_),
    .A2(net87),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07365_ (.I(_01773_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07366_ (.A1(_01765_),
    .A2(_01770_),
    .A3(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07367_ (.I(_01775_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07368_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07369_ (.I(_01771_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07370_ (.I(_01778_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07371_ (.I(net87),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07372_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07373_ (.I(_00500_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07374_ (.A1(_01782_),
    .A2(_00756_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07375_ (.A1(\as2650.cycle[6] ),
    .A2(_00549_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07376_ (.A1(\as2650.addr_buff[7] ),
    .A2(_00608_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07377_ (.A1(_00598_),
    .A2(_01019_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07378_ (.A1(_01785_),
    .A2(_01786_),
    .B(_00992_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07379_ (.A1(_00841_),
    .A2(_01784_),
    .B1(_01787_),
    .B2(_00519_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07380_ (.A1(_05734_),
    .A2(_00985_),
    .A3(_05823_),
    .A4(_00641_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07381_ (.A1(_00515_),
    .A2(_00992_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07382_ (.A1(_00986_),
    .A2(_00714_),
    .A3(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07383_ (.A1(_01011_),
    .A2(_01788_),
    .A3(_01789_),
    .B1(_01791_),
    .B2(_00609_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07384_ (.A1(_00972_),
    .A2(_01792_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07385_ (.A1(_00927_),
    .A2(_00933_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07386_ (.A1(_00952_),
    .A2(_01794_),
    .A3(_01102_),
    .B(_01763_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07387_ (.I(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07388_ (.A1(_05696_),
    .A2(_01783_),
    .B(_01793_),
    .C(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07389_ (.I(_01797_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07390_ (.I(net59),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07391_ (.A1(_01799_),
    .A2(_01768_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07392_ (.I(_01800_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07393_ (.I(_01801_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07394_ (.I(_01802_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07395_ (.I(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07396_ (.I(_01804_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07397_ (.A1(_01779_),
    .A2(_01781_),
    .A3(_01798_),
    .A4(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07398_ (.I(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07399_ (.A1(\as2650.stack[13][0] ),
    .A2(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07400_ (.A1(_00500_),
    .A2(_00756_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07401_ (.A1(_01793_),
    .A2(_01796_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07402_ (.A1(_00666_),
    .A2(_01809_),
    .B(_01810_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07403_ (.I(_01811_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07404_ (.I(net89),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07405_ (.A1(_01767_),
    .A2(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07406_ (.I(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07407_ (.A1(_01774_),
    .A2(_01812_),
    .A3(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07408_ (.I(_01816_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07409_ (.I(net93),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07410_ (.I(_01818_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07411_ (.I(_01819_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07412_ (.I(_01796_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07413_ (.I(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07414_ (.A1(_01100_),
    .A2(_01821_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07415_ (.A1(_01820_),
    .A2(_01822_),
    .B(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07416_ (.I(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07417_ (.I(_01775_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07418_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07419_ (.A1(_01817_),
    .A2(_01825_),
    .B(_01827_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07420_ (.A1(_01761_),
    .A2(_01777_),
    .B1(_01808_),
    .B2(_01828_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07421_ (.I(net86),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07422_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07423_ (.I(_01830_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07424_ (.I(_01831_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07425_ (.I(_01816_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07426_ (.I(net92),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07427_ (.I(_01834_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07428_ (.I(_01835_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07429_ (.A1(_01239_),
    .A2(_01822_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07430_ (.A1(_01836_),
    .A2(_01822_),
    .B(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07431_ (.I(_01838_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_01806_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07433_ (.A1(\as2650.stack[13][1] ),
    .A2(_01840_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07434_ (.A1(_01833_),
    .A2(_01839_),
    .B(_01841_),
    .C(_01776_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07435_ (.A1(_01832_),
    .A2(_01777_),
    .B(_01842_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07436_ (.I(net49),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07437_ (.I(_01843_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07438_ (.I(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07439_ (.I(_01845_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07440_ (.I(_00435_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07441_ (.A1(_00640_),
    .A2(_01762_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07442_ (.A1(_01016_),
    .A2(_01848_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07443_ (.I(_01794_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07444_ (.A1(_01850_),
    .A2(_01142_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07445_ (.A1(_01849_),
    .A2(_01851_),
    .ZN(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07446_ (.I(_01852_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07447_ (.I(net57),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07448_ (.I(_01854_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07449_ (.A1(_01855_),
    .A2(_01852_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07450_ (.A1(_01847_),
    .A2(_01853_),
    .B(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07451_ (.I(_01857_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07452_ (.A1(\as2650.stack[13][2] ),
    .A2(_01840_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07453_ (.A1(_01833_),
    .A2(_01858_),
    .B(_01859_),
    .C(_01826_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07454_ (.A1(_01846_),
    .A2(_01777_),
    .B(_01860_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07455_ (.I(_01068_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07456_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07457_ (.I(_01862_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(\as2650.stack[13][3] ),
    .A2(_01807_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07459_ (.I(_01852_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07460_ (.I(net58),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07461_ (.I(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07462_ (.A1(_01867_),
    .A2(_01853_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07463_ (.A1(_01354_),
    .A2(_01865_),
    .B(_01868_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07464_ (.I(_01869_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07465_ (.I(_01826_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07466_ (.A1(_01817_),
    .A2(_01870_),
    .B(_01871_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07467_ (.A1(_01863_),
    .A2(_01777_),
    .B1(_01864_),
    .B2(_01872_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07468_ (.I(_01459_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07469_ (.I(_01873_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07470_ (.I(_01776_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07471_ (.I(_01816_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07472_ (.I(_01876_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07473_ (.I(net60),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07474_ (.I(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07475_ (.I(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07476_ (.I(_01821_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07477_ (.A1(_01419_),
    .A2(_01821_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07478_ (.A1(_01880_),
    .A2(_01881_),
    .B(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07479_ (.I(_01883_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07480_ (.A1(_01877_),
    .A2(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07481_ (.A1(\as2650.stack[13][4] ),
    .A2(_01840_),
    .B(_01871_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07482_ (.A1(_01874_),
    .A2(_01875_),
    .B1(_01885_),
    .B2(_01886_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07483_ (.I(net52),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07484_ (.I(_01887_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07485_ (.I(_01888_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07486_ (.I(_01889_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07487_ (.A1(\as2650.stack[13][5] ),
    .A2(_01807_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07488_ (.I(net61),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07489_ (.I(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07490_ (.I(_01893_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07491_ (.I(_01822_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07492_ (.I(_01496_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07493_ (.A1(_01896_),
    .A2(_01881_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07494_ (.A1(_01894_),
    .A2(_01895_),
    .B(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07495_ (.I(_01898_),
    .Z(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07496_ (.A1(_01817_),
    .A2(_01899_),
    .B(_01871_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07497_ (.A1(_01890_),
    .A2(_01875_),
    .B1(_01891_),
    .B2(_01900_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07498_ (.I(_05705_),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07499_ (.I(_01901_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07500_ (.I(_01902_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(\as2650.stack[13][6] ),
    .A2(_01807_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07502_ (.I(net62),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07503_ (.I(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _07504_ (.I(_01906_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07505_ (.I(_01583_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07506_ (.A1(_01908_),
    .A2(_01881_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07507_ (.A1(_01907_),
    .A2(_01895_),
    .B(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07508_ (.I(_01910_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07509_ (.A1(_01817_),
    .A2(_01911_),
    .B(_01871_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07510_ (.A1(_01903_),
    .A2(_01875_),
    .B1(_01904_),
    .B2(_01912_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07511_ (.I(_05717_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07512_ (.I(_01913_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\as2650.stack[13][7] ),
    .A2(_01840_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07514_ (.I(_01677_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07515_ (.I(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07516_ (.I(net63),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07517_ (.I(_01918_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07518_ (.A1(_01919_),
    .A2(_01853_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07519_ (.A1(_01917_),
    .A2(_01853_),
    .B(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07520_ (.I(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07521_ (.A1(_01833_),
    .A2(_01922_),
    .B(_01776_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07522_ (.A1(_01914_),
    .A2(_01875_),
    .B1(_01915_),
    .B2(_01923_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07523_ (.I(\as2650.r123[0][0] ),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07524_ (.I(_00927_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07525_ (.A1(_01925_),
    .A2(_00928_),
    .A3(_00686_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07526_ (.I(_01926_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07527_ (.I(_01927_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07528_ (.A1(_00936_),
    .A2(_01928_),
    .B(_01142_),
    .C(_01141_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07529_ (.I(_01925_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07530_ (.I(_00928_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07531_ (.I(_01931_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _07532_ (.A1(_01930_),
    .A2(_01932_),
    .A3(_01029_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07533_ (.A1(_00513_),
    .A2(_01929_),
    .A3(_01933_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07534_ (.I(_01934_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07535_ (.I(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07536_ (.I(_01136_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07537_ (.I(_01933_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07538_ (.I(_00934_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07539_ (.I(_01939_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07540_ (.A1(_01141_),
    .A2(_01940_),
    .A3(_01142_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07541_ (.I(_01941_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07542_ (.I(_01942_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07543_ (.A1(net59),
    .A2(net89),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07544_ (.I(_01944_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07545_ (.I(net87),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07546_ (.A1(_01771_),
    .A2(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07547_ (.A1(_01945_),
    .A2(_01947_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07548_ (.A1(_01771_),
    .A2(_01769_),
    .B(_01946_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07549_ (.A1(_01948_),
    .A2(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07550_ (.I(_01950_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07551_ (.I(_01951_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07552_ (.I(_01952_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07553_ (.A1(net70),
    .A2(_01944_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07554_ (.I(_01954_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07555_ (.I(_01955_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07556_ (.I(_01956_),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07557_ (.A1(_01767_),
    .A2(net48),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07558_ (.I(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07559_ (.I(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07560_ (.I(_01960_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07561_ (.I(_01961_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07562_ (.I(_01944_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07563_ (.I(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07564_ (.I(_01964_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07565_ (.I(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07566_ (.A1(_01766_),
    .A2(_01768_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07567_ (.I(_01967_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07568_ (.I(_01968_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07569_ (.I(_01969_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07570_ (.A1(\as2650.stack[7][8] ),
    .A2(_01966_),
    .B1(_01970_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07571_ (.I(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07572_ (.A1(\as2650.stack[4][8] ),
    .A2(_01804_),
    .B1(_01962_),
    .B2(\as2650.stack[5][8] ),
    .C(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07573_ (.I(_01945_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07574_ (.I(_01974_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07575_ (.I(_01975_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07576_ (.I(_01800_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07577_ (.I(_01977_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07578_ (.I(_01978_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07579_ (.I(_01959_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07580_ (.I(_01980_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07581_ (.I(_01981_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07582_ (.A1(\as2650.stack[3][8] ),
    .A2(_01976_),
    .B1(_01979_),
    .B2(\as2650.stack[0][8] ),
    .C1(_01982_),
    .C2(\as2650.stack[1][8] ),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07583_ (.I(_01968_),
    .Z(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07584_ (.I(_01984_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07585_ (.I(_01985_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07586_ (.I(_01954_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07587_ (.I(_01987_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07588_ (.I(_01988_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07589_ (.A1(\as2650.stack[2][8] ),
    .A2(_01986_),
    .B(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07590_ (.A1(_01957_),
    .A2(_01973_),
    .B1(_01983_),
    .B2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07591_ (.I(_01974_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07592_ (.I(_01992_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07593_ (.A1(\as2650.stack[11][8] ),
    .A2(_01993_),
    .B1(_01979_),
    .B2(\as2650.stack[8][8] ),
    .C1(\as2650.stack[9][8] ),
    .C2(_01982_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07594_ (.I(_01970_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07595_ (.I(_01987_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07596_ (.I(_01996_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07597_ (.A1(\as2650.stack[10][8] ),
    .A2(_01995_),
    .B(_01997_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07598_ (.I(_01996_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07599_ (.I(_01958_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07600_ (.I(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07601_ (.I(_02001_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07602_ (.A1(\as2650.stack[15][8] ),
    .A2(_01966_),
    .B1(_02002_),
    .B2(\as2650.stack[13][8] ),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07603_ (.I(_01801_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07604_ (.I(_02004_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07605_ (.A1(\as2650.stack[12][8] ),
    .A2(_02005_),
    .B1(_01985_),
    .B2(\as2650.stack[14][8] ),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07606_ (.A1(_01999_),
    .A2(_02003_),
    .A3(_02006_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07607_ (.I(_01950_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07608_ (.I(_02008_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07609_ (.A1(_01994_),
    .A2(_01998_),
    .B(_02007_),
    .C(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07610_ (.A1(_01953_),
    .A2(_01991_),
    .B(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07611_ (.A1(_01143_),
    .A2(_01929_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07612_ (.I(_02012_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07613_ (.I(_01941_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07614_ (.A1(_01138_),
    .A2(_02014_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07615_ (.A1(_01943_),
    .A2(_02011_),
    .B(_02013_),
    .C(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07616_ (.A1(_01937_),
    .A2(_01938_),
    .B(_01935_),
    .C(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07617_ (.A1(_01924_),
    .A2(_01936_),
    .B(_02017_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07618_ (.I(\as2650.r123[0][1] ),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07619_ (.I(_01232_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07620_ (.I(_01950_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07621_ (.I(_02020_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07622_ (.I(_02021_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07623_ (.I(_01961_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07624_ (.A1(\as2650.stack[7][9] ),
    .A2(_01975_),
    .B1(_01970_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07625_ (.I(_02024_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07626_ (.A1(\as2650.stack[4][9] ),
    .A2(_01979_),
    .B1(_02023_),
    .B2(\as2650.stack[5][9] ),
    .C(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07627_ (.A1(\as2650.stack[3][9] ),
    .A2(_01976_),
    .B1(_01979_),
    .B2(\as2650.stack[0][9] ),
    .C1(_01982_),
    .C2(\as2650.stack[1][9] ),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07628_ (.A1(\as2650.stack[2][9] ),
    .A2(_01995_),
    .B(_01997_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07629_ (.A1(_01957_),
    .A2(_02026_),
    .B1(_02027_),
    .B2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07630_ (.I(net70),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07631_ (.A1(_02030_),
    .A2(_01963_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07632_ (.I(_02031_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07633_ (.I(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07634_ (.I(_02005_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07635_ (.I(_02002_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07636_ (.A1(\as2650.stack[8][9] ),
    .A2(_02034_),
    .B1(_02035_),
    .B2(\as2650.stack[9][9] ),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07637_ (.I(_01966_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07638_ (.A1(\as2650.stack[11][9] ),
    .A2(_02037_),
    .B1(_01986_),
    .B2(\as2650.stack[10][9] ),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07639_ (.A1(_02033_),
    .A2(_02036_),
    .A3(_02038_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07640_ (.I(_01963_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07641_ (.I(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07642_ (.I(_02041_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07643_ (.I(_01800_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07644_ (.I(_02043_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07645_ (.I(_02044_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07646_ (.A1(\as2650.stack[15][9] ),
    .A2(_02042_),
    .B1(_02045_),
    .B2(\as2650.stack[12][9] ),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07647_ (.I(_01967_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07648_ (.I(_02047_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07649_ (.I(_02048_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07650_ (.I(_02049_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07651_ (.I(_02000_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_02051_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07653_ (.A1(\as2650.stack[14][9] ),
    .A2(_02050_),
    .B1(_02052_),
    .B2(\as2650.stack[13][9] ),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07654_ (.A1(_01999_),
    .A2(_02046_),
    .A3(_02053_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07655_ (.A1(_02009_),
    .A2(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07656_ (.A1(_02022_),
    .A2(_02029_),
    .B1(_02039_),
    .B2(_02055_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07657_ (.A1(_01240_),
    .A2(_02014_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07658_ (.I(_02012_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07659_ (.A1(_01943_),
    .A2(_02056_),
    .B(_02057_),
    .C(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07660_ (.A1(_02019_),
    .A2(_01938_),
    .B(_01935_),
    .C(_02059_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07661_ (.A1(_02018_),
    .A2(_01936_),
    .B(_02060_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07662_ (.I(\as2650.r123[0][2] ),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07663_ (.I(_01301_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07664_ (.I(_01934_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07665_ (.I(_02009_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07666_ (.I(_01989_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07667_ (.I(_02045_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07668_ (.I(_02051_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07669_ (.I(_02067_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07670_ (.I(_02041_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07671_ (.I(_02047_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07672_ (.I(_02070_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07673_ (.I(_02071_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07674_ (.A1(\as2650.stack[7][10] ),
    .A2(_02069_),
    .B1(_02072_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07675_ (.I(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07676_ (.A1(\as2650.stack[4][10] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\as2650.stack[5][10] ),
    .C(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07677_ (.I(_02049_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07678_ (.I(_02076_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07679_ (.A1(\as2650.stack[0][10] ),
    .A2(_02066_),
    .B1(_02077_),
    .B2(\as2650.stack[2][10] ),
    .C1(\as2650.stack[1][10] ),
    .C2(_02068_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07680_ (.I(_01993_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07681_ (.A1(\as2650.stack[3][10] ),
    .A2(_02079_),
    .B(_01957_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07682_ (.A1(_02065_),
    .A2(_02075_),
    .B1(_02078_),
    .B2(_02080_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07683_ (.I(_02033_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07684_ (.I(_02044_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07685_ (.I(_02083_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07686_ (.I(_02052_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07687_ (.A1(\as2650.stack[8][10] ),
    .A2(_02084_),
    .B1(_02085_),
    .B2(\as2650.stack[9][10] ),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07688_ (.I(_02072_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07689_ (.A1(\as2650.stack[11][10] ),
    .A2(_02079_),
    .B1(_02087_),
    .B2(\as2650.stack[10][10] ),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07690_ (.A1(_02082_),
    .A2(_02086_),
    .A3(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07691_ (.I(_01956_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07692_ (.I(_01975_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07693_ (.A1(\as2650.stack[15][10] ),
    .A2(_02091_),
    .B1(_02035_),
    .B2(\as2650.stack[13][10] ),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07694_ (.A1(\as2650.stack[12][10] ),
    .A2(_01804_),
    .B1(_01986_),
    .B2(\as2650.stack[14][10] ),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07695_ (.A1(_02090_),
    .A2(_02092_),
    .A3(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07696_ (.A1(_01953_),
    .A2(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07697_ (.A1(_02064_),
    .A2(_02081_),
    .B1(_02089_),
    .B2(_02095_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07698_ (.A1(_01247_),
    .A2(_02014_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07699_ (.A1(_01943_),
    .A2(_02096_),
    .B(_02097_),
    .C(_02058_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07700_ (.A1(_02062_),
    .A2(_01938_),
    .B(_02063_),
    .C(_02098_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07701_ (.A1(_02061_),
    .A2(_01936_),
    .B(_02099_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07702_ (.I(\as2650.r123[0][3] ),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07703_ (.I(_01370_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07704_ (.I(_01941_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07705_ (.I(_02045_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07706_ (.I(_02067_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07707_ (.I(_01964_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07708_ (.I(_02105_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07709_ (.A1(\as2650.stack[7][11] ),
    .A2(_02106_),
    .B1(_02076_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07710_ (.I(_02107_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07711_ (.A1(\as2650.stack[4][11] ),
    .A2(_02103_),
    .B1(_02104_),
    .B2(\as2650.stack[5][11] ),
    .C(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07712_ (.I(_02004_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07713_ (.I(_02110_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07714_ (.I(_01985_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07715_ (.I(_02001_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07716_ (.I(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07717_ (.A1(\as2650.stack[0][11] ),
    .A2(_02111_),
    .B1(_02112_),
    .B2(\as2650.stack[2][11] ),
    .C1(\as2650.stack[1][11] ),
    .C2(_02114_),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07718_ (.I(_02069_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07719_ (.A1(\as2650.stack[3][11] ),
    .A2(_02116_),
    .B(_02090_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07720_ (.A1(_02065_),
    .A2(_02109_),
    .B1(_02115_),
    .B2(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07721_ (.I(_02083_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07722_ (.I(_02052_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07723_ (.A1(\as2650.stack[8][11] ),
    .A2(_02119_),
    .B1(_02120_),
    .B2(\as2650.stack[9][11] ),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07724_ (.I(_02072_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07725_ (.A1(\as2650.stack[11][11] ),
    .A2(_02116_),
    .B1(_02122_),
    .B2(\as2650.stack[10][11] ),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07726_ (.A1(_02082_),
    .A2(_02121_),
    .A3(_02123_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07727_ (.I(_01956_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07728_ (.A1(\as2650.stack[15][11] ),
    .A2(_01976_),
    .B1(_02023_),
    .B2(\as2650.stack[13][11] ),
    .ZN(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07729_ (.I(_01803_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07730_ (.A1(\as2650.stack[12][11] ),
    .A2(_02127_),
    .B1(_01995_),
    .B2(\as2650.stack[14][11] ),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07731_ (.A1(_02125_),
    .A2(_02126_),
    .A3(_02128_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07732_ (.A1(_02022_),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07733_ (.A1(_02064_),
    .A2(_02118_),
    .B1(_02124_),
    .B2(_02130_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07734_ (.I(_01323_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07735_ (.I(_02132_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07736_ (.A1(_02133_),
    .A2(_02014_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07737_ (.A1(_02102_),
    .A2(_02131_),
    .B(_02134_),
    .C(_02058_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07738_ (.A1(_02101_),
    .A2(_01938_),
    .B(_02063_),
    .C(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07739_ (.A1(_02100_),
    .A2(_01936_),
    .B(_02136_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07740_ (.I(_01935_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07741_ (.I(_01933_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07742_ (.A1(\as2650.stack[7][12] ),
    .A2(_02106_),
    .B1(_02076_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07743_ (.I(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07744_ (.A1(\as2650.stack[4][12] ),
    .A2(_02103_),
    .B1(_02104_),
    .B2(\as2650.stack[5][12] ),
    .C(_02140_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07745_ (.A1(\as2650.stack[0][12] ),
    .A2(_02034_),
    .B1(_02112_),
    .B2(\as2650.stack[2][12] ),
    .C1(\as2650.stack[1][12] ),
    .C2(_02114_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07746_ (.I(_02106_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07747_ (.A1(\as2650.stack[3][12] ),
    .A2(_02143_),
    .B(_02125_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07748_ (.A1(_01957_),
    .A2(_02141_),
    .B1(_02142_),
    .B2(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07749_ (.A1(\as2650.stack[8][12] ),
    .A2(_02119_),
    .B1(_02120_),
    .B2(\as2650.stack[9][12] ),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07750_ (.A1(\as2650.stack[11][12] ),
    .A2(_02116_),
    .B1(_02122_),
    .B2(\as2650.stack[10][12] ),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07751_ (.A1(_02033_),
    .A2(_02146_),
    .A3(_02147_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07752_ (.A1(\as2650.stack[15][12] ),
    .A2(_01976_),
    .B1(_02127_),
    .B2(\as2650.stack[12][12] ),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07753_ (.I(_02070_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07754_ (.I(_02150_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07755_ (.A1(\as2650.stack[14][12] ),
    .A2(_02151_),
    .B1(_02023_),
    .B2(\as2650.stack[13][12] ),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07756_ (.A1(_01989_),
    .A2(_02149_),
    .A3(_02152_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07757_ (.A1(_02022_),
    .A2(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07758_ (.A1(_01953_),
    .A2(_02145_),
    .B1(_02148_),
    .B2(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07759_ (.I(_01419_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07760_ (.A1(_02156_),
    .A2(_01942_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07761_ (.A1(_02102_),
    .A2(_02155_),
    .B(_02157_),
    .C(_02013_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07762_ (.A1(_01457_),
    .A2(_02138_),
    .B(_02063_),
    .C(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07763_ (.A1(_01464_),
    .A2(_02137_),
    .B(_02159_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07764_ (.I(_01536_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07765_ (.A1(\as2650.stack[7][13] ),
    .A2(_02042_),
    .B1(_02050_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07766_ (.I(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07767_ (.A1(\as2650.stack[4][13] ),
    .A2(_02103_),
    .B1(_02068_),
    .B2(\as2650.stack[5][13] ),
    .C(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07768_ (.A1(\as2650.stack[3][13] ),
    .A2(_02037_),
    .B1(_02111_),
    .B2(\as2650.stack[0][13] ),
    .C1(_02114_),
    .C2(\as2650.stack[1][13] ),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07769_ (.I(_02072_),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07770_ (.A1(\as2650.stack[2][13] ),
    .A2(_02165_),
    .B(_02090_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07771_ (.A1(_02065_),
    .A2(_02163_),
    .B1(_02164_),
    .B2(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07772_ (.A1(\as2650.stack[8][13] ),
    .A2(_02119_),
    .B1(_02120_),
    .B2(\as2650.stack[9][13] ),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07773_ (.I(_02069_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07774_ (.A1(\as2650.stack[11][13] ),
    .A2(_02169_),
    .B1(_02122_),
    .B2(\as2650.stack[10][13] ),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07775_ (.A1(_02082_),
    .A2(_02168_),
    .A3(_02170_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07776_ (.A1(\as2650.stack[15][13] ),
    .A2(_02091_),
    .B1(_02127_),
    .B2(\as2650.stack[12][13] ),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07777_ (.A1(\as2650.stack[14][13] ),
    .A2(_01995_),
    .B1(_01962_),
    .B2(\as2650.stack[13][13] ),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07778_ (.A1(_02125_),
    .A2(_02172_),
    .A3(_02173_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07779_ (.A1(_02022_),
    .A2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07780_ (.A1(_02064_),
    .A2(_02167_),
    .B1(_02171_),
    .B2(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07781_ (.A1(_01896_),
    .A2(_01942_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07782_ (.A1(_02102_),
    .A2(_02176_),
    .B(_02177_),
    .C(_02013_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07783_ (.A1(_02160_),
    .A2(_02138_),
    .B(_02063_),
    .C(_02178_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07784_ (.A1(_01542_),
    .A2(_02137_),
    .B(_02179_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07785_ (.I(_01624_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07786_ (.A1(\as2650.stack[7][14] ),
    .A2(_02042_),
    .B1(_02050_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07787_ (.I(_02181_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07788_ (.A1(\as2650.stack[4][14] ),
    .A2(_02066_),
    .B1(_02068_),
    .B2(\as2650.stack[5][14] ),
    .C(_02182_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07789_ (.A1(\as2650.stack[0][14] ),
    .A2(_02111_),
    .B1(_02077_),
    .B2(\as2650.stack[2][14] ),
    .C1(\as2650.stack[1][14] ),
    .C2(_02104_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07790_ (.A1(\as2650.stack[3][14] ),
    .A2(_02169_),
    .B(_02090_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07791_ (.A1(_02065_),
    .A2(_02183_),
    .B1(_02184_),
    .B2(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07792_ (.A1(\as2650.stack[8][14] ),
    .A2(_02111_),
    .B1(_02077_),
    .B2(\as2650.stack[10][14] ),
    .C1(_02114_),
    .C2(\as2650.stack[9][14] ),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07793_ (.A1(\as2650.stack[11][14] ),
    .A2(_02143_),
    .B(_02125_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07794_ (.A1(\as2650.stack[15][14] ),
    .A2(_01993_),
    .B1(_02052_),
    .B2(\as2650.stack[13][14] ),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07795_ (.A1(\as2650.stack[12][14] ),
    .A2(_02083_),
    .B1(_02151_),
    .B2(\as2650.stack[14][14] ),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07796_ (.A1(_01989_),
    .A2(_02189_),
    .A3(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _07797_ (.A1(_02187_),
    .A2(_02188_),
    .B(_02191_),
    .C(_02009_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07798_ (.A1(_02064_),
    .A2(_02186_),
    .B(_02192_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07799_ (.A1(_01908_),
    .A2(_01942_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07800_ (.A1(_02102_),
    .A2(_02193_),
    .B(_02194_),
    .C(_02013_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07801_ (.A1(_02180_),
    .A2(_02138_),
    .B(_01934_),
    .C(_02195_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07802_ (.A1(_01645_),
    .A2(_02137_),
    .B(_02196_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07803_ (.I(\as2650.r123[0][7] ),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07804_ (.I(_01718_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07805_ (.I(_01917_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07806_ (.A1(_02199_),
    .A2(_01943_),
    .A3(_02058_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07807_ (.A1(_02198_),
    .A2(_02138_),
    .B(_01934_),
    .C(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07808_ (.A1(_02197_),
    .A2(_02137_),
    .B(_02201_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07809_ (.I(_01799_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07810_ (.I(_01768_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07811_ (.A1(_02202_),
    .A2(_02203_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07812_ (.I(_02204_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07813_ (.A1(_01774_),
    .A2(_01812_),
    .A3(_02205_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07814_ (.I(_02206_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07815_ (.I(_02207_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07816_ (.I(_01851_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07817_ (.I(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07818_ (.I(_01852_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07819_ (.I(net91),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07820_ (.I(_02212_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07821_ (.I(_02213_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07822_ (.A1(_01151_),
    .A2(_02210_),
    .B1(_02211_),
    .B2(_02214_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07823_ (.I(_02215_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07824_ (.I(_01764_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07825_ (.I(_01773_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07826_ (.I(_01814_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07827_ (.A1(_02217_),
    .A2(_02218_),
    .A3(_02219_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07829_ (.I(_02221_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07830_ (.I(_02206_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07831_ (.A1(\as2650.stack[14][8] ),
    .A2(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07832_ (.A1(_02208_),
    .A2(_02216_),
    .B(_02222_),
    .C(_02224_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07833_ (.I(net65),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07834_ (.I(_02225_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07835_ (.A1(_01237_),
    .A2(_02210_),
    .B1(_02211_),
    .B2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07836_ (.I(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07837_ (.I(_02206_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07838_ (.A1(\as2650.stack[14][9] ),
    .A2(_02229_),
    .ZN(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07839_ (.I(_02221_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07840_ (.A1(_02208_),
    .A2(_02228_),
    .B(_02230_),
    .C(_02231_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07841_ (.I(net66),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07842_ (.I(_02232_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07843_ (.I(_02233_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07844_ (.A1(_01313_),
    .A2(_02210_),
    .B1(_02211_),
    .B2(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07845_ (.I(_02235_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07846_ (.A1(\as2650.stack[14][10] ),
    .A2(_02229_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07847_ (.A1(_02208_),
    .A2(_02236_),
    .B(_02237_),
    .C(_02231_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07848_ (.I(net67),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07849_ (.I(_02238_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07850_ (.I(_02239_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07851_ (.A1(_01385_),
    .A2(_02210_),
    .B1(_02211_),
    .B2(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07852_ (.I(_02241_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07853_ (.A1(\as2650.stack[14][11] ),
    .A2(_02229_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07854_ (.A1(_02208_),
    .A2(_02242_),
    .B(_02243_),
    .C(_02231_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07855_ (.I(_02207_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07856_ (.I(net68),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _07857_ (.I(_02245_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07858_ (.A1(_01634_),
    .A2(_02209_),
    .B1(_01865_),
    .B2(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07859_ (.I(_02247_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07860_ (.A1(\as2650.stack[14][12] ),
    .A2(_02229_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07861_ (.A1(_02244_),
    .A2(_02248_),
    .B(_02249_),
    .C(_02231_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07862_ (.I(net69),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07863_ (.A1(_01631_),
    .A2(_02209_),
    .B1(_01865_),
    .B2(_02250_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07864_ (.I(_02251_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07865_ (.A1(\as2650.stack[14][13] ),
    .A2(_02207_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07866_ (.A1(_02244_),
    .A2(_02252_),
    .B(_02253_),
    .C(_02222_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07867_ (.I(_01647_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07868_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07869_ (.I(_02255_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07870_ (.A1(_02256_),
    .A2(_02209_),
    .B1(_01865_),
    .B2(net90),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07871_ (.I(_02257_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07872_ (.A1(\as2650.stack[14][14] ),
    .A2(_02207_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07873_ (.A1(_02244_),
    .A2(_02258_),
    .B(_02259_),
    .C(_02222_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07874_ (.I(_01876_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07875_ (.A1(\as2650.stack[13][8] ),
    .A2(_01833_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07876_ (.I(_01826_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07877_ (.A1(_02260_),
    .A2(_02216_),
    .B(_02261_),
    .C(_02262_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07878_ (.I(_01816_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07879_ (.A1(\as2650.stack[13][9] ),
    .A2(_02263_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07880_ (.A1(_02260_),
    .A2(_02228_),
    .B(_02264_),
    .C(_02262_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07881_ (.A1(\as2650.stack[13][10] ),
    .A2(_02263_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07882_ (.A1(_02260_),
    .A2(_02236_),
    .B(_02265_),
    .C(_02262_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07883_ (.A1(\as2650.stack[13][11] ),
    .A2(_02263_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07884_ (.A1(_02260_),
    .A2(_02242_),
    .B(_02266_),
    .C(_02262_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07885_ (.A1(\as2650.stack[13][12] ),
    .A2(_02263_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07886_ (.A1(_01877_),
    .A2(_02248_),
    .B(_02267_),
    .C(_01827_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07887_ (.A1(\as2650.stack[13][13] ),
    .A2(_01876_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07888_ (.A1(_01877_),
    .A2(_02252_),
    .B(_02268_),
    .C(_01827_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07889_ (.A1(\as2650.stack[13][14] ),
    .A2(_01876_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07890_ (.A1(_01877_),
    .A2(_02258_),
    .B(_02269_),
    .C(_01827_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07891_ (.A1(_02030_),
    .A2(net73),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07892_ (.I(_02270_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07893_ (.A1(_02217_),
    .A2(_02219_),
    .A3(_02271_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07894_ (.I(_02272_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07895_ (.I(_02273_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07896_ (.I(_01798_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07897_ (.I(_02120_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07898_ (.I(_01947_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07899_ (.A1(_02275_),
    .A2(_02276_),
    .A3(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07900_ (.I(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07901_ (.A1(\as2650.stack[10][0] ),
    .A2(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07902_ (.I(_01824_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07903_ (.I(_02281_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07904_ (.I(_01811_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07905_ (.A1(_02283_),
    .A2(_02205_),
    .A3(_02271_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07906_ (.I(_02284_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07907_ (.I(_02272_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07908_ (.I(_02286_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07909_ (.A1(_02282_),
    .A2(_02285_),
    .B(_02287_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07910_ (.A1(_01761_),
    .A2(_02274_),
    .B1(_02280_),
    .B2(_02288_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07911_ (.I(_01830_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(\as2650.stack[10][1] ),
    .A2(_02279_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07913_ (.I(_01839_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07914_ (.I(_02286_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07915_ (.A1(_02291_),
    .A2(_02285_),
    .B(_02292_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07916_ (.A1(_02289_),
    .A2(_02274_),
    .B1(_02290_),
    .B2(_02293_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(\as2650.stack[10][2] ),
    .A2(_02279_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07918_ (.I(_01857_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07919_ (.I(_02284_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07920_ (.A1(_02295_),
    .A2(_02296_),
    .B(_02292_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07921_ (.A1(_01846_),
    .A2(_02274_),
    .B1(_02294_),
    .B2(_02297_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07922_ (.I(_01869_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07923_ (.I(_02284_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07924_ (.I(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(_02298_),
    .A2(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07926_ (.I(_02278_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07927_ (.A1(\as2650.stack[10][3] ),
    .A2(_02302_),
    .B(_02292_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07928_ (.A1(_01863_),
    .A2(_02274_),
    .B1(_02301_),
    .B2(_02303_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07929_ (.I(_02286_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07930_ (.A1(\as2650.stack[10][4] ),
    .A2(_02279_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07931_ (.A1(_01884_),
    .A2(_02296_),
    .B(_02292_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07932_ (.A1(_01874_),
    .A2(_02304_),
    .B1(_02305_),
    .B2(_02306_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07933_ (.I(_01898_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07934_ (.A1(_02307_),
    .A2(_02285_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07935_ (.A1(\as2650.stack[10][5] ),
    .A2(_02302_),
    .B(_02273_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07936_ (.A1(_01890_),
    .A2(_02304_),
    .B1(_02308_),
    .B2(_02309_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07937_ (.I(_01910_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07938_ (.A1(_02310_),
    .A2(_02285_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07939_ (.A1(\as2650.stack[10][6] ),
    .A2(_02302_),
    .B(_02273_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07940_ (.A1(_01903_),
    .A2(_02304_),
    .B1(_02311_),
    .B2(_02312_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07941_ (.A1(\as2650.stack[10][7] ),
    .A2(_02302_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07942_ (.I(_01921_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07943_ (.A1(_02314_),
    .A2(_02296_),
    .B(_02273_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07944_ (.A1(_01914_),
    .A2(_02304_),
    .B1(_02313_),
    .B2(_02315_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07945_ (.A1(_01769_),
    .A2(_02218_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07946_ (.A1(_02316_),
    .A2(_01797_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07947_ (.I(_02317_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07948_ (.I(_02318_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07949_ (.I(_02317_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07950_ (.A1(\as2650.stack[12][8] ),
    .A2(_02320_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07951_ (.I(_01799_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07952_ (.A1(_02322_),
    .A2(_01813_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07953_ (.I(_02323_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07954_ (.A1(_02217_),
    .A2(_02324_),
    .A3(_02270_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07955_ (.I(_02325_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07956_ (.I(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07957_ (.A1(_02216_),
    .A2(_02319_),
    .B(_02321_),
    .C(_02327_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07958_ (.I(_02318_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07959_ (.A1(\as2650.stack[12][9] ),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07960_ (.A1(_02228_),
    .A2(_02319_),
    .B(_02327_),
    .C(_02329_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07961_ (.A1(\as2650.stack[12][10] ),
    .A2(_02328_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07962_ (.A1(_02236_),
    .A2(_02319_),
    .B(_02327_),
    .C(_02330_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07963_ (.A1(\as2650.stack[12][11] ),
    .A2(_02328_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07964_ (.A1(_02242_),
    .A2(_02319_),
    .B(_02327_),
    .C(_02331_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07965_ (.I(_02318_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07966_ (.I(_02326_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07967_ (.A1(\as2650.stack[12][12] ),
    .A2(_02320_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07968_ (.A1(_02248_),
    .A2(_02332_),
    .B(_02333_),
    .C(_02334_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07969_ (.A1(\as2650.stack[12][13] ),
    .A2(_02320_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07970_ (.A1(_02252_),
    .A2(_02332_),
    .B(_02333_),
    .C(_02335_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07971_ (.A1(\as2650.stack[12][14] ),
    .A2(_02320_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07972_ (.A1(_02258_),
    .A2(_02332_),
    .B(_02333_),
    .C(_02336_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07973_ (.I(_02324_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07974_ (.A1(_02283_),
    .A2(_02337_),
    .A3(_02271_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07975_ (.I(_02338_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07976_ (.I(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07977_ (.A1(\as2650.stack[11][8] ),
    .A2(_02339_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07978_ (.I(_01764_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07979_ (.I(_02204_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07980_ (.A1(_02342_),
    .A2(_02343_),
    .A3(_02270_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07981_ (.I(_02344_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07982_ (.I(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07983_ (.A1(_02216_),
    .A2(_02340_),
    .B(_02341_),
    .C(_02346_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07984_ (.I(_02338_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07985_ (.A1(\as2650.stack[11][9] ),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07986_ (.A1(_02228_),
    .A2(_02340_),
    .B(_02346_),
    .C(_02348_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07987_ (.I(_02338_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07988_ (.A1(\as2650.stack[11][10] ),
    .A2(_02349_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07989_ (.A1(_02236_),
    .A2(_02340_),
    .B(_02346_),
    .C(_02350_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07990_ (.A1(\as2650.stack[11][11] ),
    .A2(_02349_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07991_ (.A1(_02242_),
    .A2(_02340_),
    .B(_02346_),
    .C(_02351_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07992_ (.I(_02339_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07993_ (.I(_02345_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07994_ (.A1(\as2650.stack[11][12] ),
    .A2(_02349_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07995_ (.A1(_02248_),
    .A2(_02352_),
    .B(_02353_),
    .C(_02354_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07996_ (.A1(\as2650.stack[11][13] ),
    .A2(_02349_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07997_ (.A1(_02252_),
    .A2(_02352_),
    .B(_02353_),
    .C(_02355_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07998_ (.A1(\as2650.stack[11][14] ),
    .A2(_02339_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07999_ (.A1(_02258_),
    .A2(_02352_),
    .B(_02353_),
    .C(_02356_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08000_ (.I(_00890_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08001_ (.A1(_00937_),
    .A2(_00686_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08002_ (.A1(_02357_),
    .A2(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08003_ (.A1(_01925_),
    .A2(_00568_),
    .A3(_00470_),
    .A4(_01337_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08004_ (.A1(_00998_),
    .A2(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08005_ (.A1(_02359_),
    .A2(_02361_),
    .B(_00766_),
    .C(_00837_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08006_ (.I(_02362_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _08007_ (.I(_00892_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08008_ (.A1(_01916_),
    .A2(_02364_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08009_ (.A1(_01932_),
    .A2(_00554_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08010_ (.A1(_00836_),
    .A2(net77),
    .B(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08011_ (.A1(_00938_),
    .A2(_02365_),
    .B1(_02367_),
    .B2(_02361_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08012_ (.A1(_00763_),
    .A2(_00603_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08013_ (.I(_02369_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08014_ (.A1(net4),
    .A2(_02363_),
    .B1(_02368_),
    .B2(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08015_ (.A1(_00755_),
    .A2(_02371_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08016_ (.I(_01760_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08017_ (.I(_02220_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08018_ (.I(_02373_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08019_ (.I(_01962_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08020_ (.A1(_01779_),
    .A2(_01781_),
    .A3(_01798_),
    .A4(_02375_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08021_ (.I(_02376_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08022_ (.A1(\as2650.stack[14][0] ),
    .A2(_02377_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08023_ (.A1(_01825_),
    .A2(_02223_),
    .B(_02373_),
    .C(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08024_ (.A1(_02372_),
    .A2(_02374_),
    .B(_02379_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08025_ (.I(_01838_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08026_ (.A1(\as2650.stack[14][1] ),
    .A2(_02377_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08027_ (.A1(_02380_),
    .A2(_02223_),
    .B(_02221_),
    .C(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08028_ (.A1(_01832_),
    .A2(_02374_),
    .B(_02382_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08029_ (.I(_02376_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08030_ (.A1(\as2650.stack[14][2] ),
    .A2(_02383_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08031_ (.I(_02206_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08032_ (.A1(_02295_),
    .A2(_02385_),
    .B(_02222_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08033_ (.A1(_01846_),
    .A2(_02374_),
    .B1(_02384_),
    .B2(_02386_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08034_ (.A1(\as2650.stack[14][3] ),
    .A2(_02383_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08035_ (.I(_01869_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08036_ (.I(_02221_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08037_ (.A1(_02388_),
    .A2(_02385_),
    .B(_02389_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08038_ (.A1(_01863_),
    .A2(_02374_),
    .B1(_02387_),
    .B2(_02390_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08039_ (.I(_02373_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08040_ (.I(_01883_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08041_ (.I(_02392_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08042_ (.A1(_02393_),
    .A2(_02244_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08043_ (.A1(\as2650.stack[14][4] ),
    .A2(_02377_),
    .B(_02389_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08044_ (.A1(_01874_),
    .A2(_02391_),
    .B1(_02394_),
    .B2(_02395_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08045_ (.A1(_02307_),
    .A2(_02385_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08046_ (.A1(\as2650.stack[14][5] ),
    .A2(_02377_),
    .B(_02389_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08047_ (.A1(_01890_),
    .A2(_02391_),
    .B1(_02396_),
    .B2(_02397_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08048_ (.I(_01901_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08049_ (.A1(\as2650.stack[14][6] ),
    .A2(_02383_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08050_ (.A1(_02310_),
    .A2(_02385_),
    .B(_02389_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08051_ (.A1(_02398_),
    .A2(_02391_),
    .B1(_02399_),
    .B2(_02400_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08052_ (.A1(\as2650.stack[14][7] ),
    .A2(_02383_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08053_ (.I(_01921_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08054_ (.A1(_02402_),
    .A2(_02223_),
    .B(_02373_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08055_ (.A1(_01914_),
    .A2(_02391_),
    .B1(_02401_),
    .B2(_02403_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08056_ (.I(_02215_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08057_ (.I(_02299_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08058_ (.A1(\as2650.stack[10][8] ),
    .A2(_02296_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08059_ (.I(_02286_),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08060_ (.A1(_02404_),
    .A2(_02405_),
    .B(_02406_),
    .C(_02407_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08061_ (.I(_02227_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08062_ (.I(_02284_),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08063_ (.A1(\as2650.stack[10][9] ),
    .A2(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08064_ (.A1(_02408_),
    .A2(_02405_),
    .B(_02410_),
    .C(_02407_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08065_ (.I(_02235_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08066_ (.A1(\as2650.stack[10][10] ),
    .A2(_02409_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08067_ (.A1(_02411_),
    .A2(_02405_),
    .B(_02412_),
    .C(_02407_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08068_ (.I(_02241_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08069_ (.A1(\as2650.stack[10][11] ),
    .A2(_02409_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08070_ (.A1(_02413_),
    .A2(_02405_),
    .B(_02414_),
    .C(_02407_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08071_ (.I(_02247_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08072_ (.A1(\as2650.stack[10][12] ),
    .A2(_02409_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08073_ (.A1(_02415_),
    .A2(_02300_),
    .B(_02416_),
    .C(_02287_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08074_ (.I(_02251_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08075_ (.A1(\as2650.stack[10][13] ),
    .A2(_02299_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08076_ (.A1(_02417_),
    .A2(_02300_),
    .B(_02418_),
    .C(_02287_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08077_ (.I(_02257_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08078_ (.A1(\as2650.stack[10][14] ),
    .A2(_02299_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08079_ (.A1(_02419_),
    .A2(_02300_),
    .B(_02420_),
    .C(_02287_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08080_ (.A1(_02217_),
    .A2(_02218_),
    .A3(_02337_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08081_ (.I(_02421_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08082_ (.I(_02422_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08083_ (.I(_02169_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08084_ (.I(_01797_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08085_ (.A1(_01779_),
    .A2(_01780_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08086_ (.I(_02426_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08087_ (.A1(_02424_),
    .A2(_02425_),
    .A3(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08088_ (.I(_02428_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(\as2650.stack[0][0] ),
    .A2(_02429_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08090_ (.I(_01812_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08091_ (.A1(_02116_),
    .A2(_02426_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08092_ (.A1(_02431_),
    .A2(_02432_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08093_ (.I(_02433_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08094_ (.I(_02421_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08095_ (.I(_02435_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08096_ (.A1(_02282_),
    .A2(_02434_),
    .B(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08097_ (.A1(_01761_),
    .A2(_02423_),
    .B1(_02430_),
    .B2(_02437_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08098_ (.A1(\as2650.stack[0][1] ),
    .A2(_02429_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08099_ (.I(_02435_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08100_ (.A1(_02291_),
    .A2(_02434_),
    .B(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08101_ (.A1(_02289_),
    .A2(_02423_),
    .B1(_02438_),
    .B2(_02440_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08102_ (.I(_01844_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(\as2650.stack[0][2] ),
    .A2(_02429_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08104_ (.A1(_02295_),
    .A2(_02434_),
    .B(_02439_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08105_ (.A1(_02441_),
    .A2(_02423_),
    .B1(_02442_),
    .B2(_02443_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08106_ (.I(_01862_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08107_ (.I(_02433_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08108_ (.I(_02445_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(_02298_),
    .A2(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08110_ (.I(_02428_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08111_ (.A1(\as2650.stack[0][3] ),
    .A2(_02448_),
    .B(_02439_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08112_ (.A1(_02444_),
    .A2(_02423_),
    .B1(_02447_),
    .B2(_02449_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08113_ (.I(_02435_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(_02393_),
    .A2(_02434_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08115_ (.A1(\as2650.stack[0][4] ),
    .A2(_02448_),
    .B(_02439_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08116_ (.A1(_01874_),
    .A2(_02450_),
    .B1(_02451_),
    .B2(_02452_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08117_ (.I(_01888_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08118_ (.A1(\as2650.stack[0][5] ),
    .A2(_02429_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08119_ (.I(_02433_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08120_ (.A1(_02307_),
    .A2(_02455_),
    .B(_02422_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08121_ (.A1(_02453_),
    .A2(_02450_),
    .B1(_02454_),
    .B2(_02456_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08122_ (.A1(\as2650.stack[0][6] ),
    .A2(_02448_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08123_ (.A1(_02310_),
    .A2(_02455_),
    .B(_02422_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08124_ (.A1(_02398_),
    .A2(_02450_),
    .B1(_02457_),
    .B2(_02458_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08125_ (.I(_01913_),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08126_ (.A1(\as2650.stack[0][7] ),
    .A2(_02448_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08127_ (.A1(_02402_),
    .A2(_02455_),
    .B(_02422_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08128_ (.A1(_02459_),
    .A2(_02450_),
    .B1(_02460_),
    .B2(_02461_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08129_ (.I(_02445_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08130_ (.A1(\as2650.stack[0][8] ),
    .A2(_02455_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08131_ (.I(_02435_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08132_ (.A1(_02404_),
    .A2(_02462_),
    .B(_02463_),
    .C(_02464_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08133_ (.I(_02433_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08134_ (.A1(\as2650.stack[0][9] ),
    .A2(_02465_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08135_ (.A1(_02408_),
    .A2(_02462_),
    .B(_02466_),
    .C(_02464_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08136_ (.A1(\as2650.stack[0][10] ),
    .A2(_02465_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08137_ (.A1(_02411_),
    .A2(_02462_),
    .B(_02467_),
    .C(_02464_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08138_ (.A1(\as2650.stack[0][11] ),
    .A2(_02465_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08139_ (.A1(_02413_),
    .A2(_02462_),
    .B(_02468_),
    .C(_02464_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08140_ (.A1(\as2650.stack[0][12] ),
    .A2(_02465_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08141_ (.A1(_02415_),
    .A2(_02446_),
    .B(_02469_),
    .C(_02436_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08142_ (.A1(\as2650.stack[0][13] ),
    .A2(_02445_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08143_ (.A1(_02417_),
    .A2(_02446_),
    .B(_02470_),
    .C(_02436_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08144_ (.A1(\as2650.stack[0][14] ),
    .A2(_02445_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08145_ (.A1(_02419_),
    .A2(_02446_),
    .B(_02471_),
    .C(_02436_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08146_ (.A1(_02431_),
    .A2(_01948_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08148_ (.I(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08149_ (.A1(\as2650.stack[8][8] ),
    .A2(_02473_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08150_ (.I(_01764_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08151_ (.I(_01946_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_01772_),
    .A2(_02477_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08153_ (.I(_02478_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08154_ (.A1(_02476_),
    .A2(_02324_),
    .A3(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08155_ (.I(_02480_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08156_ (.I(_02481_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08157_ (.A1(_02404_),
    .A2(_02474_),
    .B(_02475_),
    .C(_02482_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08158_ (.I(_02472_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08159_ (.A1(\as2650.stack[8][9] ),
    .A2(_02483_),
    .ZN(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08160_ (.A1(_02408_),
    .A2(_02474_),
    .B(_02482_),
    .C(_02484_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08161_ (.I(_02472_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08162_ (.A1(\as2650.stack[8][10] ),
    .A2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08163_ (.A1(_02411_),
    .A2(_02474_),
    .B(_02482_),
    .C(_02486_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08164_ (.A1(\as2650.stack[8][11] ),
    .A2(_02485_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08165_ (.A1(_02413_),
    .A2(_02474_),
    .B(_02482_),
    .C(_02487_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08166_ (.I(_02473_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08167_ (.I(_02481_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08168_ (.A1(\as2650.stack[8][12] ),
    .A2(_02485_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08169_ (.A1(_02415_),
    .A2(_02488_),
    .B(_02489_),
    .C(_02490_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08170_ (.A1(\as2650.stack[8][13] ),
    .A2(_02485_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08171_ (.A1(_02417_),
    .A2(_02488_),
    .B(_02489_),
    .C(_02491_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08172_ (.A1(\as2650.stack[8][14] ),
    .A2(_02473_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08173_ (.A1(_02419_),
    .A2(_02488_),
    .B(_02489_),
    .C(_02492_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08174_ (.I(_02478_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08175_ (.A1(_02283_),
    .A2(_02337_),
    .A3(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08176_ (.I(_02494_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08177_ (.I(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08178_ (.A1(\as2650.stack[7][8] ),
    .A2(_02495_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08179_ (.A1(_02342_),
    .A2(_02343_),
    .A3(_02493_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08180_ (.I(_02498_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08181_ (.I(_02499_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08182_ (.A1(_02404_),
    .A2(_02496_),
    .B(_02497_),
    .C(_02500_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08183_ (.I(_02494_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08184_ (.A1(\as2650.stack[7][9] ),
    .A2(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08185_ (.A1(_02408_),
    .A2(_02496_),
    .B(_02500_),
    .C(_02502_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08186_ (.I(_02494_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08187_ (.A1(\as2650.stack[7][10] ),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08188_ (.A1(_02411_),
    .A2(_02496_),
    .B(_02500_),
    .C(_02504_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08189_ (.A1(\as2650.stack[7][11] ),
    .A2(_02503_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08190_ (.A1(_02413_),
    .A2(_02496_),
    .B(_02500_),
    .C(_02505_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08191_ (.I(_02495_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08192_ (.I(_02499_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08193_ (.A1(\as2650.stack[7][12] ),
    .A2(_02503_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08194_ (.A1(_02415_),
    .A2(_02506_),
    .B(_02507_),
    .C(_02508_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08195_ (.A1(\as2650.stack[7][13] ),
    .A2(_02503_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08196_ (.A1(_02417_),
    .A2(_02506_),
    .B(_02507_),
    .C(_02509_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08197_ (.A1(\as2650.stack[7][14] ),
    .A2(_02495_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08198_ (.A1(_02419_),
    .A2(_02506_),
    .B(_02507_),
    .C(_02510_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08199_ (.I(_01004_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08200_ (.I(_02511_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08201_ (.A1(_00636_),
    .A2(_02512_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08202_ (.I(_00763_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08203_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08204_ (.A1(_02515_),
    .A2(_00873_),
    .B(_00703_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _08205_ (.A1(_05728_),
    .A2(_00506_),
    .A3(_02513_),
    .B(_02516_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08206_ (.A1(_00704_),
    .A2(_00756_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08207_ (.A1(_00502_),
    .A2(_05704_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(_02519_),
    .A2(_02369_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08209_ (.I(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08210_ (.A1(_00631_),
    .A2(_00695_),
    .A3(_01189_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08211_ (.I(_00906_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08212_ (.A1(_00789_),
    .A2(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08213_ (.A1(_01460_),
    .A2(_02370_),
    .A3(_02524_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08214_ (.A1(_02521_),
    .A2(_02522_),
    .B(_02525_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08215_ (.A1(_00478_),
    .A2(_00687_),
    .A3(_00956_),
    .A4(_01004_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08216_ (.A1(_02517_),
    .A2(_02518_),
    .A3(_02526_),
    .A4(_02527_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08217_ (.A1(_00773_),
    .A2(_00890_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08218_ (.A1(_00934_),
    .A2(_01926_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08219_ (.A1(_00696_),
    .A2(_02529_),
    .A3(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08220_ (.A1(_00929_),
    .A2(_00811_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08221_ (.A1(_00948_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08222_ (.A1(_02533_),
    .A2(_00949_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08223_ (.A1(_01850_),
    .A2(_00938_),
    .A3(_02531_),
    .A4(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08224_ (.A1(_00884_),
    .A2(_00888_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08225_ (.A1(_00630_),
    .A2(_00695_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08226_ (.A1(_00891_),
    .A2(_02537_),
    .A3(_02521_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08227_ (.A1(_00568_),
    .A2(_01337_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08228_ (.A1(_00955_),
    .A2(_00697_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08229_ (.A1(_02539_),
    .A2(_02540_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08230_ (.A1(_00537_),
    .A2(_02360_),
    .A3(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08231_ (.A1(_02536_),
    .A2(_02538_),
    .A3(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08232_ (.A1(_00763_),
    .A2(_00535_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08233_ (.I(_02544_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08234_ (.I(_02541_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08235_ (.A1(_00705_),
    .A2(_00780_),
    .A3(_02545_),
    .A4(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08236_ (.A1(_00887_),
    .A2(_00625_),
    .B(_02521_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08237_ (.A1(_00764_),
    .A2(_00505_),
    .A3(_00509_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08238_ (.A1(_02548_),
    .A2(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08239_ (.A1(_02535_),
    .A2(_02543_),
    .A3(_02547_),
    .A4(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08240_ (.A1(_00952_),
    .A2(_00496_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08241_ (.A1(_00946_),
    .A2(_02552_),
    .A3(_00949_),
    .A4(_02511_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08242_ (.A1(_00689_),
    .A2(_01004_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08243_ (.A1(_01112_),
    .A2(_00930_),
    .A3(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08244_ (.A1(_02553_),
    .A2(_02555_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08245_ (.A1(_00782_),
    .A2(_01206_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08246_ (.A1(_02514_),
    .A2(_00873_),
    .A3(_00500_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08247_ (.I(_02558_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08248_ (.I(_02559_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08249_ (.A1(_00891_),
    .A2(_00631_),
    .A3(_02521_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08250_ (.I(_00527_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08251_ (.A1(_05728_),
    .A2(_00878_),
    .A3(_02512_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08252_ (.A1(_01279_),
    .A2(_00837_),
    .A3(_02562_),
    .A4(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08253_ (.A1(_02557_),
    .A2(_02560_),
    .B(_02561_),
    .C(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08254_ (.A1(_00466_),
    .A2(_02523_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08255_ (.A1(_00923_),
    .A2(_01926_),
    .A3(_02566_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08256_ (.A1(_02520_),
    .A2(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08257_ (.I(_02357_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08258_ (.I(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08259_ (.I(_02570_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08260_ (.A1(_01925_),
    .A2(_00922_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08261_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08262_ (.I(_02573_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08263_ (.A1(_00773_),
    .A2(_02571_),
    .A3(_00691_),
    .A4(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08264_ (.A1(_02556_),
    .A2(_02565_),
    .A3(_02568_),
    .A4(_02575_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08265_ (.A1(_02528_),
    .A2(_02551_),
    .A3(_02576_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08266_ (.I(_00632_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08267_ (.I(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08268_ (.I(_02364_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08269_ (.I(_02580_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _08270_ (.I(_01500_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08271_ (.I(_02582_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08272_ (.I(_02583_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _08273_ (.A1(_01931_),
    .A2(_02360_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08274_ (.I(_00892_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08275_ (.I(_02586_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08276_ (.I(_02587_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08277_ (.I(_02570_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08278_ (.I(_01500_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08279_ (.I(_02590_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08280_ (.A1(_02589_),
    .A2(_02591_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08281_ (.I(net75),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08282_ (.A1(_01896_),
    .A2(_02588_),
    .B1(_02592_),
    .B2(_02593_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08283_ (.A1(_02581_),
    .A2(_02584_),
    .A3(_02585_),
    .B(_02594_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08284_ (.I(_01782_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08285_ (.I(_02596_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08286_ (.I(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08287_ (.A1(_02579_),
    .A2(_02595_),
    .B(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08288_ (.A1(_02593_),
    .A2(_02577_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08289_ (.A1(_02577_),
    .A2(_02599_),
    .B(_02600_),
    .C(_00830_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08290_ (.I(_02215_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08291_ (.A1(_01812_),
    .A2(_02343_),
    .A3(_02479_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08292_ (.I(_02602_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08293_ (.I(_02603_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08294_ (.I(_02604_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08295_ (.A1(\as2650.stack[6][8] ),
    .A2(_02604_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08296_ (.A1(_02476_),
    .A2(_02219_),
    .A3(_02479_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08297_ (.I(_02607_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08298_ (.I(_02608_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08299_ (.A1(_02601_),
    .A2(_02605_),
    .B(_02606_),
    .C(_02609_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08300_ (.I(_02227_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08301_ (.I(_02603_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08302_ (.A1(\as2650.stack[6][9] ),
    .A2(_02611_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08303_ (.A1(_02610_),
    .A2(_02605_),
    .B(_02609_),
    .C(_02612_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08304_ (.I(_02235_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08305_ (.I(_02608_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08306_ (.I(_02603_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08307_ (.A1(\as2650.stack[6][10] ),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08308_ (.A1(_02613_),
    .A2(_02605_),
    .B(_02614_),
    .C(_02616_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08309_ (.I(_02241_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08310_ (.A1(\as2650.stack[6][11] ),
    .A2(_02615_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08311_ (.A1(_02617_),
    .A2(_02605_),
    .B(_02614_),
    .C(_02618_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08312_ (.I(_02247_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08313_ (.I(_02602_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08314_ (.I(_02620_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08315_ (.A1(\as2650.stack[6][12] ),
    .A2(_02615_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08316_ (.A1(_02619_),
    .A2(_02621_),
    .B(_02614_),
    .C(_02622_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08317_ (.I(_02251_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08318_ (.A1(\as2650.stack[6][13] ),
    .A2(_02615_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08319_ (.A1(_02623_),
    .A2(_02621_),
    .B(_02614_),
    .C(_02624_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08320_ (.I(_02257_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08321_ (.I(_02607_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08322_ (.A1(\as2650.stack[6][14] ),
    .A2(_02604_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08323_ (.A1(_02625_),
    .A2(_02621_),
    .B(_02626_),
    .C(_02627_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08324_ (.I(_01811_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08325_ (.A1(_02628_),
    .A2(_01815_),
    .A3(_02493_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08326_ (.I(_02629_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08327_ (.I(_02630_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08328_ (.A1(\as2650.stack[5][8] ),
    .A2(_02630_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08329_ (.A1(_02342_),
    .A2(_01770_),
    .A3(_02479_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08330_ (.I(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08331_ (.I(_02634_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08332_ (.A1(_02601_),
    .A2(_02631_),
    .B(_02632_),
    .C(_02635_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08333_ (.I(_02629_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08334_ (.A1(\as2650.stack[5][9] ),
    .A2(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08335_ (.A1(_02610_),
    .A2(_02631_),
    .B(_02635_),
    .C(_02637_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08336_ (.I(_02629_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08337_ (.A1(\as2650.stack[5][10] ),
    .A2(_02638_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08338_ (.A1(_02613_),
    .A2(_02631_),
    .B(_02635_),
    .C(_02639_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08339_ (.A1(\as2650.stack[5][11] ),
    .A2(_02638_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08340_ (.A1(_02617_),
    .A2(_02631_),
    .B(_02635_),
    .C(_02640_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08341_ (.I(_02630_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08342_ (.I(_02634_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08343_ (.A1(\as2650.stack[5][12] ),
    .A2(_02638_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08344_ (.A1(_02619_),
    .A2(_02641_),
    .B(_02642_),
    .C(_02643_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08345_ (.A1(\as2650.stack[5][13] ),
    .A2(_02638_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08346_ (.A1(_02623_),
    .A2(_02641_),
    .B(_02642_),
    .C(_02644_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08347_ (.A1(\as2650.stack[5][14] ),
    .A2(_02630_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08348_ (.A1(_02625_),
    .A2(_02641_),
    .B(_02642_),
    .C(_02645_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08349_ (.A1(_01770_),
    .A2(_02431_),
    .A3(_02493_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08350_ (.I(_02646_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08351_ (.I(_02647_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08352_ (.A1(\as2650.stack[4][8] ),
    .A2(_02647_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08353_ (.A1(_02165_),
    .A2(_02426_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08354_ (.A1(_01765_),
    .A2(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08355_ (.I(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08356_ (.I(_02652_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08357_ (.A1(_02601_),
    .A2(_02648_),
    .B(_02649_),
    .C(_02653_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08358_ (.I(_02646_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08359_ (.A1(\as2650.stack[4][9] ),
    .A2(_02654_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08360_ (.A1(_02610_),
    .A2(_02648_),
    .B(_02653_),
    .C(_02655_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08361_ (.A1(\as2650.stack[4][10] ),
    .A2(_02654_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08362_ (.A1(_02613_),
    .A2(_02648_),
    .B(_02653_),
    .C(_02656_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08363_ (.I(_02652_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08364_ (.A1(\as2650.stack[4][11] ),
    .A2(_02654_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08365_ (.A1(_02617_),
    .A2(_02648_),
    .B(_02657_),
    .C(_02658_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08366_ (.I(_02647_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08367_ (.A1(\as2650.stack[4][12] ),
    .A2(_02654_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08368_ (.A1(_02619_),
    .A2(_02659_),
    .B(_02657_),
    .C(_02660_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08369_ (.I(_02646_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08370_ (.A1(\as2650.stack[4][13] ),
    .A2(_02661_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08371_ (.A1(_02623_),
    .A2(_02659_),
    .B(_02657_),
    .C(_02662_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08372_ (.A1(\as2650.stack[4][14] ),
    .A2(_02661_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08373_ (.A1(_02625_),
    .A2(_02659_),
    .B(_02657_),
    .C(_02663_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08374_ (.I(_02325_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08375_ (.I(_02664_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08376_ (.I(_01797_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08377_ (.A1(_02316_),
    .A2(_02666_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08378_ (.I(_02667_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08379_ (.I(_01881_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08380_ (.I(_01819_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08381_ (.I(_02670_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08382_ (.A1(_02671_),
    .A2(_01895_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08383_ (.A1(_01138_),
    .A2(_02669_),
    .B(_02672_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08384_ (.A1(_02673_),
    .A2(_02667_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08385_ (.A1(\as2650.stack[12][0] ),
    .A2(_02668_),
    .B(_02664_),
    .C(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08386_ (.A1(_02372_),
    .A2(_02665_),
    .B(_02675_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08387_ (.I(_01239_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08388_ (.A1(_01836_),
    .A2(_01895_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08389_ (.A1(_02676_),
    .A2(_02669_),
    .B(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08390_ (.A1(_02678_),
    .A2(_02667_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08391_ (.A1(\as2650.stack[12][1] ),
    .A2(_02668_),
    .B(_02326_),
    .C(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08392_ (.A1(_01832_),
    .A2(_02665_),
    .B(_02680_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08393_ (.I(_02667_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08394_ (.A1(\as2650.stack[12][2] ),
    .A2(_02681_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08395_ (.I(_02318_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08396_ (.A1(_02295_),
    .A2(_02683_),
    .B(_02333_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08397_ (.A1(_02441_),
    .A2(_02665_),
    .B1(_02682_),
    .B2(_02684_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08398_ (.A1(_02298_),
    .A2(_02332_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08399_ (.I(_02326_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08400_ (.A1(\as2650.stack[12][3] ),
    .A2(_02668_),
    .B(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08401_ (.A1(_02444_),
    .A2(_02665_),
    .B1(_02685_),
    .B2(_02687_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08402_ (.I(_01459_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08403_ (.I(_02664_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08404_ (.A1(\as2650.stack[12][4] ),
    .A2(_02681_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08405_ (.A1(_02392_),
    .A2(_02683_),
    .B(_02686_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08406_ (.A1(_02688_),
    .A2(_02689_),
    .B1(_02690_),
    .B2(_02691_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08407_ (.A1(\as2650.stack[12][5] ),
    .A2(_02681_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08408_ (.A1(_02307_),
    .A2(_02683_),
    .B(_02686_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08409_ (.A1(_02453_),
    .A2(_02689_),
    .B1(_02692_),
    .B2(_02693_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(\as2650.stack[12][6] ),
    .A2(_02681_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08411_ (.I(_01910_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08412_ (.A1(_02695_),
    .A2(_02683_),
    .B(_02686_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08413_ (.A1(_02398_),
    .A2(_02689_),
    .B1(_02694_),
    .B2(_02696_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08414_ (.A1(\as2650.stack[12][7] ),
    .A2(_02668_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08415_ (.A1(_02402_),
    .A2(_02328_),
    .B(_02664_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08416_ (.A1(_02459_),
    .A2(_02689_),
    .B1(_02697_),
    .B2(_02698_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08417_ (.A1(_02431_),
    .A2(_02650_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08418_ (.I(_02699_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08419_ (.I(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08420_ (.A1(\as2650.stack[3][8] ),
    .A2(_02700_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08421_ (.I(_02030_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08422_ (.A1(_02703_),
    .A2(_02477_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08423_ (.A1(_02342_),
    .A2(_02343_),
    .A3(_02704_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08424_ (.I(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08425_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08426_ (.A1(_02601_),
    .A2(_02701_),
    .B(_02702_),
    .C(_02707_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08427_ (.I(_02699_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08428_ (.A1(\as2650.stack[3][9] ),
    .A2(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08429_ (.A1(_02610_),
    .A2(_02701_),
    .B(_02707_),
    .C(_02709_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08430_ (.I(_02699_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08431_ (.A1(\as2650.stack[3][10] ),
    .A2(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08432_ (.A1(_02613_),
    .A2(_02701_),
    .B(_02707_),
    .C(_02711_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08433_ (.A1(\as2650.stack[3][11] ),
    .A2(_02710_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08434_ (.A1(_02617_),
    .A2(_02701_),
    .B(_02707_),
    .C(_02712_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08435_ (.I(_02700_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08436_ (.I(_02706_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08437_ (.A1(\as2650.stack[3][12] ),
    .A2(_02710_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08438_ (.A1(_02619_),
    .A2(_02713_),
    .B(_02714_),
    .C(_02715_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08439_ (.A1(\as2650.stack[3][13] ),
    .A2(_02710_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08440_ (.A1(_02623_),
    .A2(_02713_),
    .B(_02714_),
    .C(_02716_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08441_ (.A1(\as2650.stack[3][14] ),
    .A2(_02700_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08442_ (.A1(_02625_),
    .A2(_02713_),
    .B(_02714_),
    .C(_02717_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08443_ (.I(_02215_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08444_ (.A1(_02628_),
    .A2(_02205_),
    .A3(_02704_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08445_ (.I(_02719_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08446_ (.I(_02720_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08447_ (.A1(\as2650.stack[2][8] ),
    .A2(_02720_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08448_ (.A1(_02476_),
    .A2(_02219_),
    .A3(_02704_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08449_ (.I(_02723_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08450_ (.I(_02724_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08451_ (.A1(_02718_),
    .A2(_02721_),
    .B(_02722_),
    .C(_02725_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08452_ (.I(_02227_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08453_ (.I(_02719_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08454_ (.A1(\as2650.stack[2][9] ),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08455_ (.A1(_02726_),
    .A2(_02721_),
    .B(_02725_),
    .C(_02728_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08456_ (.I(_02235_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08457_ (.I(_02719_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08458_ (.A1(\as2650.stack[2][10] ),
    .A2(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08459_ (.A1(_02729_),
    .A2(_02721_),
    .B(_02725_),
    .C(_02731_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08460_ (.I(_02241_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08461_ (.A1(\as2650.stack[2][11] ),
    .A2(_02730_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08462_ (.A1(_02732_),
    .A2(_02721_),
    .B(_02725_),
    .C(_02733_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08463_ (.I(_02247_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08464_ (.I(_02720_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08465_ (.I(_02724_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08466_ (.A1(\as2650.stack[2][12] ),
    .A2(_02730_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08467_ (.A1(_02734_),
    .A2(_02735_),
    .B(_02736_),
    .C(_02737_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08468_ (.I(_02251_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08469_ (.A1(\as2650.stack[2][13] ),
    .A2(_02730_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08470_ (.A1(_02738_),
    .A2(_02735_),
    .B(_02736_),
    .C(_02739_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08471_ (.I(_02257_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08472_ (.A1(\as2650.stack[2][14] ),
    .A2(_02720_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08473_ (.A1(_02740_),
    .A2(_02735_),
    .B(_02736_),
    .C(_02741_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08474_ (.A1(_02628_),
    .A2(_01815_),
    .A3(_02704_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08475_ (.I(_02742_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08476_ (.I(_02743_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08477_ (.A1(\as2650.stack[1][8] ),
    .A2(_02743_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08478_ (.A1(_01765_),
    .A2(_02432_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08479_ (.I(_02746_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08480_ (.I(_02747_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08481_ (.A1(_02718_),
    .A2(_02744_),
    .B(_02745_),
    .C(_02748_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08482_ (.I(_02742_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08483_ (.A1(\as2650.stack[1][9] ),
    .A2(_02749_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08484_ (.A1(_02726_),
    .A2(_02744_),
    .B(_02748_),
    .C(_02750_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08485_ (.I(_02742_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08486_ (.A1(\as2650.stack[1][10] ),
    .A2(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08487_ (.A1(_02729_),
    .A2(_02744_),
    .B(_02748_),
    .C(_02752_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08488_ (.A1(\as2650.stack[1][11] ),
    .A2(_02751_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08489_ (.A1(_02732_),
    .A2(_02744_),
    .B(_02748_),
    .C(_02753_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08490_ (.I(_02743_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08491_ (.I(_02747_),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08492_ (.A1(\as2650.stack[1][12] ),
    .A2(_02751_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08493_ (.A1(_02734_),
    .A2(_02754_),
    .B(_02755_),
    .C(_02756_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08494_ (.A1(\as2650.stack[1][13] ),
    .A2(_02751_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08495_ (.A1(_02738_),
    .A2(_02754_),
    .B(_02755_),
    .C(_02757_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08496_ (.A1(\as2650.stack[1][14] ),
    .A2(_02743_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08497_ (.A1(_02740_),
    .A2(_02754_),
    .B(_02755_),
    .C(_02758_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08498_ (.A1(_01774_),
    .A2(_02283_),
    .A3(_02337_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08499_ (.I(_02759_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08500_ (.I(_02760_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08501_ (.A1(\as2650.stack[15][8] ),
    .A2(_02760_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08502_ (.A1(_02476_),
    .A2(_02218_),
    .A3(_02205_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08503_ (.I(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08504_ (.I(_02764_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08505_ (.A1(_02718_),
    .A2(_02761_),
    .B(_02762_),
    .C(_02765_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08506_ (.I(_02759_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08507_ (.A1(\as2650.stack[15][9] ),
    .A2(_02766_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08508_ (.A1(_02726_),
    .A2(_02761_),
    .B(_02765_),
    .C(_02767_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08509_ (.I(_02759_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08510_ (.A1(\as2650.stack[15][10] ),
    .A2(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08511_ (.A1(_02729_),
    .A2(_02761_),
    .B(_02765_),
    .C(_02769_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08512_ (.A1(\as2650.stack[15][11] ),
    .A2(_02768_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08513_ (.A1(_02732_),
    .A2(_02761_),
    .B(_02765_),
    .C(_02770_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08514_ (.I(_02760_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08515_ (.I(_02764_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08516_ (.A1(\as2650.stack[15][12] ),
    .A2(_02768_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08517_ (.A1(_02734_),
    .A2(_02771_),
    .B(_02772_),
    .C(_02773_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08518_ (.A1(\as2650.stack[15][13] ),
    .A2(_02768_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08519_ (.A1(_02738_),
    .A2(_02771_),
    .B(_02772_),
    .C(_02774_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08520_ (.A1(\as2650.stack[15][14] ),
    .A2(_02760_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08521_ (.A1(_02740_),
    .A2(_02771_),
    .B(_02772_),
    .C(_02775_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08522_ (.A1(_00782_),
    .A2(_00814_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08523_ (.I(_02566_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08524_ (.A1(_00898_),
    .A2(_02776_),
    .B(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08525_ (.A1(_00804_),
    .A2(_00886_),
    .A3(_00529_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08526_ (.A1(_05718_),
    .A2(_00803_),
    .A3(_00917_),
    .B(_00952_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08527_ (.A1(_01848_),
    .A2(_02567_),
    .A3(_02779_),
    .A4(_02780_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08528_ (.I(_00891_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08529_ (.A1(_00824_),
    .A2(_00635_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08530_ (.A1(_00781_),
    .A2(_00536_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08531_ (.A1(_00643_),
    .A2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08532_ (.A1(_02783_),
    .A2(_02785_),
    .B(_00953_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08533_ (.A1(_02357_),
    .A2(_00644_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08534_ (.A1(_02782_),
    .A2(_00954_),
    .B(_02786_),
    .C(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08535_ (.A1(_02778_),
    .A2(_02781_),
    .A3(_02788_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08536_ (.I(_00896_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08537_ (.A1(_00536_),
    .A2(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08538_ (.A1(_00813_),
    .A2(_00820_),
    .A3(_00898_),
    .A4(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08539_ (.A1(_00735_),
    .A2(_00897_),
    .A3(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08540_ (.A1(_00640_),
    .A2(_00462_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08541_ (.A1(_00953_),
    .A2(_01931_),
    .A3(_02361_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08542_ (.A1(_02794_),
    .A2(_02795_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08543_ (.A1(_02514_),
    .A2(_00496_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08544_ (.A1(_00703_),
    .A2(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08545_ (.A1(_00529_),
    .A2(_00630_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08546_ (.A1(_00887_),
    .A2(_02799_),
    .A3(_00998_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08547_ (.I(_00693_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08548_ (.A1(_02523_),
    .A2(_01206_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08549_ (.A1(_02801_),
    .A2(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08550_ (.I(_00993_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08551_ (.A1(_00875_),
    .A2(_00677_),
    .A3(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08552_ (.A1(_02798_),
    .A2(_02800_),
    .A3(_02803_),
    .A4(_02805_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08553_ (.A1(_02793_),
    .A2(_02796_),
    .A3(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_02782_),
    .A2(_00957_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08555_ (.A1(_02522_),
    .A2(_02808_),
    .B(_02557_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08556_ (.I(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08557_ (.I(_02523_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08558_ (.I(_02811_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08559_ (.A1(_02812_),
    .A2(_01939_),
    .B1(_02361_),
    .B2(_05718_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08560_ (.I(_02811_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _08561_ (.A1(_02814_),
    .A2(_02790_),
    .A3(_02799_),
    .B1(_02359_),
    .B2(_00796_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08562_ (.A1(_00705_),
    .A2(_02813_),
    .B(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08563_ (.A1(_01112_),
    .A2(_00728_),
    .A3(_02537_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08564_ (.A1(_00947_),
    .A2(_02542_),
    .A3(_02817_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08565_ (.A1(_02810_),
    .A2(_02816_),
    .A3(_02818_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08566_ (.A1(_02789_),
    .A2(_02807_),
    .A3(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08567_ (.I(_02814_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08568_ (.I(_02821_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08569_ (.I(_02822_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08570_ (.A1(_01531_),
    .A2(_01520_),
    .B(_01612_),
    .C(_01444_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08571_ (.A1(_01705_),
    .A2(_02824_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08572_ (.A1(_01051_),
    .A2(_01170_),
    .A3(_01293_),
    .A4(_01329_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08573_ (.I(_00987_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08574_ (.A1(net86),
    .A2(_01706_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08575_ (.A1(_01329_),
    .A2(_01332_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08576_ (.A1(_01071_),
    .A2(_01176_),
    .B(_01281_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08577_ (.A1(_01293_),
    .A2(_01328_),
    .A3(_02830_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08578_ (.A1(_01432_),
    .A2(_02829_),
    .A3(_02831_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_01521_),
    .A2(_01524_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08580_ (.A1(_01604_),
    .A2(_02833_),
    .B(_01613_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08581_ (.A1(_01710_),
    .A2(_02834_),
    .B(_01705_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_01699_),
    .A2(_01702_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08583_ (.A1(_02832_),
    .A2(_02825_),
    .B(_02835_),
    .C(_02836_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08584_ (.A1(_02828_),
    .A2(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08585_ (.A1(_02827_),
    .A2(_02838_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08586_ (.A1(_02825_),
    .A2(_02826_),
    .B(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08587_ (.A1(_02823_),
    .A2(_02840_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08588_ (.I(_01188_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08589_ (.A1(net80),
    .A2(_02842_),
    .A3(_01534_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08590_ (.I(_01343_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08591_ (.A1(_01299_),
    .A2(_02844_),
    .A3(_01455_),
    .A4(_01622_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08592_ (.A1(_02843_),
    .A2(_02845_),
    .B(_02827_),
    .C(_01717_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08593_ (.A1(_01582_),
    .A2(_01495_),
    .A3(_01418_),
    .A4(_02132_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08594_ (.A1(_01246_),
    .A2(_01202_),
    .A3(_01099_),
    .A4(_02847_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(_01579_),
    .A2(_00821_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08596_ (.A1(_01678_),
    .A2(_00821_),
    .A3(_02848_),
    .B1(_02849_),
    .B2(_01683_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08597_ (.I(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08598_ (.I(_00667_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08599_ (.I(_02852_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08600_ (.I(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08601_ (.A1(_02841_),
    .A2(_02846_),
    .B1(_02851_),
    .B2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08602_ (.A1(_00797_),
    .A2(_00569_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08603_ (.I(_02856_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08604_ (.I(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08605_ (.I(_00887_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08606_ (.I(_02859_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08607_ (.I(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08608_ (.I(_01116_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08609_ (.I(_02862_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08610_ (.I(_02863_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08611_ (.I(_01211_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08612_ (.I(_01252_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08613_ (.I(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08614_ (.I(_02867_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08615_ (.I(_01347_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _08616_ (.I(_02869_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08617_ (.I(_02870_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08618_ (.I(_02871_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08619_ (.I(_02872_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08620_ (.A1(_02864_),
    .A2(_02865_),
    .A3(_02868_),
    .A4(_02873_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08621_ (.I(_01409_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08622_ (.I(_02875_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08623_ (.I(_01576_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08624_ (.A1(_02876_),
    .A2(_02591_),
    .A3(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08625_ (.A1(_02874_),
    .A2(_02878_),
    .B(_00554_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08626_ (.I(_00621_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08627_ (.I(_02880_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08628_ (.A1(_02881_),
    .A2(_01673_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08629_ (.I(_00429_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08630_ (.I(_01249_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08631_ (.A1(_01345_),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08632_ (.I(_01595_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08633_ (.A1(_01579_),
    .A2(_02886_),
    .A3(_01413_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08634_ (.A1(_02883_),
    .A2(_01404_),
    .A3(_02885_),
    .A4(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08635_ (.I(_02801_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08636_ (.A1(_02889_),
    .A2(_01110_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08637_ (.A1(_01588_),
    .A2(_02890_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08638_ (.I(_02889_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08639_ (.I(_02782_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08640_ (.A1(_01677_),
    .A2(_02848_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08641_ (.I0(_02894_),
    .I1(_01583_),
    .S(_02534_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08642_ (.A1(_01930_),
    .A2(_00490_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08643_ (.I(net53),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08644_ (.A1(_02897_),
    .A2(_01575_),
    .B(_02814_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08645_ (.A1(_01931_),
    .A2(_01576_),
    .B(_02896_),
    .C(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08646_ (.A1(_02893_),
    .A2(_02895_),
    .B1(_02899_),
    .B2(_02539_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_02892_),
    .A2(_02900_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08648_ (.I(_00637_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08649_ (.A1(_01670_),
    .A2(_02902_),
    .B(_02880_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08650_ (.A1(_02891_),
    .A2(_02901_),
    .A3(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08651_ (.I(_02859_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08652_ (.A1(_02882_),
    .A2(_02888_),
    .B(_02904_),
    .C(_02905_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08653_ (.A1(_02861_),
    .A2(_02879_),
    .B(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08654_ (.A1(\as2650.stack[7][6] ),
    .A2(_02105_),
    .B1(_02049_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08655_ (.I(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08656_ (.A1(\as2650.stack[4][6] ),
    .A2(_02110_),
    .B1(_02113_),
    .B2(\as2650.stack[5][6] ),
    .C(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _08657_ (.A1(\as2650.stack[0][6] ),
    .A2(_01803_),
    .B1(_01985_),
    .B2(\as2650.stack[2][6] ),
    .C1(_02002_),
    .C2(\as2650.stack[1][6] ),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08658_ (.A1(\as2650.stack[3][6] ),
    .A2(_02042_),
    .B(_01988_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08659_ (.A1(_01999_),
    .A2(_02910_),
    .B1(_02911_),
    .B2(_02912_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08660_ (.A1(\as2650.stack[8][6] ),
    .A2(_02045_),
    .B1(_02067_),
    .B2(\as2650.stack[9][6] ),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08661_ (.A1(\as2650.stack[11][6] ),
    .A2(_02069_),
    .B1(_02050_),
    .B2(\as2650.stack[10][6] ),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08662_ (.A1(_02033_),
    .A2(_02914_),
    .A3(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08663_ (.A1(\as2650.stack[15][6] ),
    .A2(_02105_),
    .B1(_02049_),
    .B2(\as2650.stack[14][6] ),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08664_ (.I(_02917_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08665_ (.A1(\as2650.stack[12][6] ),
    .A2(_02110_),
    .B1(_02113_),
    .B2(\as2650.stack[13][6] ),
    .C(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08666_ (.A1(_01997_),
    .A2(_02919_),
    .B(_02021_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _08667_ (.A1(_01952_),
    .A2(_02913_),
    .B1(_02916_),
    .B2(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08668_ (.I(_00798_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08669_ (.A1(_02858_),
    .A2(_02907_),
    .B1(_02921_),
    .B2(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08670_ (.A1(_00678_),
    .A2(_02855_),
    .B(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08671_ (.A1(_02897_),
    .A2(_02820_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08672_ (.I(_05700_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08673_ (.A1(_02820_),
    .A2(_02924_),
    .B(_02925_),
    .C(_02926_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08674_ (.A1(_02588_),
    .A2(_02839_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08675_ (.I(_01717_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08676_ (.A1(_02827_),
    .A2(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08677_ (.A1(_02199_),
    .A2(_00917_),
    .B(_02823_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08678_ (.A1(_02927_),
    .A2(_02929_),
    .B1(_02849_),
    .B2(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08679_ (.A1(_00678_),
    .A2(_02931_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08680_ (.I(_00798_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08681_ (.I(_02031_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08682_ (.I(_01959_),
    .Z(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08683_ (.A1(\as2650.stack[8][7] ),
    .A2(_01802_),
    .B1(_02935_),
    .B2(\as2650.stack[9][7] ),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08684_ (.I(_01964_),
    .Z(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08685_ (.A1(\as2650.stack[11][7] ),
    .A2(_02937_),
    .B1(_01969_),
    .B2(\as2650.stack[10][7] ),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08686_ (.A1(_02934_),
    .A2(_02936_),
    .A3(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08687_ (.I(_01954_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08688_ (.A1(\as2650.stack[15][7] ),
    .A2(_02937_),
    .B1(_01969_),
    .B2(\as2650.stack[14][7] ),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08689_ (.A1(\as2650.stack[12][7] ),
    .A2(_01802_),
    .B1(_02935_),
    .B2(\as2650.stack[13][7] ),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08690_ (.A1(_02940_),
    .A2(_02941_),
    .A3(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_02939_),
    .A2(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08692_ (.I(_01945_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08693_ (.I(_01801_),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08694_ (.A1(\as2650.stack[7][7] ),
    .A2(_02945_),
    .B1(_02946_),
    .B2(\as2650.stack[4][7] ),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08695_ (.I(_01968_),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08696_ (.A1(\as2650.stack[6][7] ),
    .A2(_02948_),
    .B1(_01960_),
    .B2(\as2650.stack[5][7] ),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08697_ (.A1(_01955_),
    .A2(_02947_),
    .A3(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08698_ (.I(_02031_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08699_ (.A1(\as2650.stack[0][7] ),
    .A2(_02946_),
    .B1(_02948_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08700_ (.A1(\as2650.stack[3][7] ),
    .A2(_02945_),
    .B1(_01960_),
    .B2(\as2650.stack[1][7] ),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08701_ (.A1(_02951_),
    .A2(_02952_),
    .A3(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08702_ (.A1(_02020_),
    .A2(_02950_),
    .A3(_02954_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08703_ (.A1(_02008_),
    .A2(_02944_),
    .B(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08704_ (.I(_02892_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08705_ (.I(_02782_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08706_ (.I(_02958_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08707_ (.I(_00550_),
    .Z(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08708_ (.I(_02960_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08709_ (.A1(_02539_),
    .A2(_02540_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08710_ (.A1(_02961_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08711_ (.A1(_00782_),
    .A2(_01074_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08712_ (.A1(_02896_),
    .A2(_02964_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08713_ (.A1(_02871_),
    .A2(_00426_),
    .B1(_01111_),
    .B2(_01210_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08714_ (.A1(_01574_),
    .A2(_01595_),
    .B1(_01204_),
    .B2(_01253_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _08715_ (.A1(_00832_),
    .A2(_01109_),
    .B1(_01424_),
    .B2(_01408_),
    .C1(_00439_),
    .C2(_01116_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08716_ (.A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08717_ (.A1(_02590_),
    .A2(_01412_),
    .B(_02965_),
    .C(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08718_ (.A1(_05717_),
    .A2(_00832_),
    .B1(_01501_),
    .B2(_01887_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _08719_ (.A1(_01069_),
    .A2(_02862_),
    .B1(_01253_),
    .B2(_01843_),
    .C1(_01861_),
    .C2(_02870_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08720_ (.A1(_01829_),
    .A2(_01210_),
    .B1(_01408_),
    .B2(_00995_),
    .C1(_01574_),
    .C2(_01901_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08721_ (.A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08722_ (.A1(_01930_),
    .A2(_02974_),
    .B(_02964_),
    .C(_00697_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _08723_ (.I(_01408_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08724_ (.I(net29),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08725_ (.A1(_02030_),
    .A2(_01253_),
    .B1(_01574_),
    .B2(_02977_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08726_ (.A1(net74),
    .A2(_02976_),
    .B1(net77),
    .B2(_00867_),
    .C(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08727_ (.I(net9),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08728_ (.I(_02980_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08729_ (.A1(_02203_),
    .A2(_02862_),
    .B1(_02870_),
    .B2(_01946_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08730_ (.A1(_02322_),
    .A2(_02981_),
    .B1(_02582_),
    .B2(_02593_),
    .C(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08731_ (.A1(_01930_),
    .A2(_00697_),
    .A3(_02964_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08732_ (.A1(_02979_),
    .A2(_02983_),
    .B(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08733_ (.A1(_00479_),
    .A2(_00490_),
    .A3(_02539_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08734_ (.A1(_02970_),
    .A2(_02975_),
    .B(_02985_),
    .C(_02986_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08735_ (.A1(_05713_),
    .A2(_00552_),
    .A3(_02986_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08736_ (.A1(_02546_),
    .A2(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08737_ (.A1(_05713_),
    .A2(_02963_),
    .B1(_02987_),
    .B2(_02989_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08738_ (.A1(_02959_),
    .A2(_02990_),
    .B(_02365_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08739_ (.A1(_02957_),
    .A2(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(_02903_),
    .A2(_02992_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08741_ (.A1(_02861_),
    .A2(_02882_),
    .A3(_02993_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08742_ (.A1(_00870_),
    .A2(_02861_),
    .B(_02994_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08743_ (.I(_02820_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08744_ (.A1(_02933_),
    .A2(_02956_),
    .B1(_02995_),
    .B2(_02858_),
    .C(_02996_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08745_ (.I(_00828_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08746_ (.I(_02998_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08747_ (.A1(_05713_),
    .A2(_02820_),
    .B(_02999_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08748_ (.A1(_02932_),
    .A2(_02997_),
    .B(_03000_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08749_ (.I(_01760_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08750_ (.I(_02763_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08751_ (.I(_03002_),
    .Z(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08752_ (.I(_02165_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08753_ (.A1(_01779_),
    .A2(_01781_),
    .A3(_02425_),
    .A4(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08754_ (.I(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08755_ (.A1(\as2650.stack[15][0] ),
    .A2(_03006_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08756_ (.I(_02759_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08757_ (.A1(_02282_),
    .A2(_03008_),
    .B(_02772_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08758_ (.A1(_03001_),
    .A2(_03003_),
    .B1(_03007_),
    .B2(_03009_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(\as2650.stack[15][1] ),
    .A2(_03006_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08760_ (.I(_02764_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08761_ (.A1(_02291_),
    .A2(_03008_),
    .B(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08762_ (.A1(_02289_),
    .A2(_03003_),
    .B1(_03010_),
    .B2(_03012_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08763_ (.A1(\as2650.stack[15][2] ),
    .A2(_03006_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08764_ (.I(_01857_),
    .Z(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08765_ (.A1(_03014_),
    .A2(_03008_),
    .B(_03011_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08766_ (.A1(_02441_),
    .A2(_03003_),
    .B1(_03013_),
    .B2(_03015_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08767_ (.A1(\as2650.stack[15][3] ),
    .A2(_03006_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08768_ (.A1(_02388_),
    .A2(_02766_),
    .B(_03011_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08769_ (.A1(_02444_),
    .A2(_03003_),
    .B1(_03016_),
    .B2(_03017_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08770_ (.I(_02764_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08771_ (.A1(_02393_),
    .A2(_02771_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08772_ (.I(_03005_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08773_ (.A1(\as2650.stack[15][4] ),
    .A2(_03020_),
    .B(_03011_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08774_ (.A1(_02688_),
    .A2(_03018_),
    .B1(_03019_),
    .B2(_03021_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08775_ (.A1(\as2650.stack[15][5] ),
    .A2(_03020_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08776_ (.I(_01898_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08777_ (.A1(_03023_),
    .A2(_02766_),
    .B(_03002_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08778_ (.A1(_02453_),
    .A2(_03018_),
    .B1(_03022_),
    .B2(_03024_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08779_ (.A1(\as2650.stack[15][6] ),
    .A2(_03020_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08780_ (.A1(_02695_),
    .A2(_02766_),
    .B(_03002_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08781_ (.A1(_02398_),
    .A2(_03018_),
    .B1(_03025_),
    .B2(_03026_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08782_ (.A1(_02314_),
    .A2(_03008_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08783_ (.A1(\as2650.stack[15][7] ),
    .A2(_03020_),
    .B(_03002_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08784_ (.A1(_02459_),
    .A2(_03018_),
    .B1(_03027_),
    .B2(_03028_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08785_ (.I(_02480_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08786_ (.I(_03029_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08787_ (.A1(_02424_),
    .A2(_02425_),
    .A3(_02277_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08788_ (.I(_03031_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08789_ (.A1(\as2650.stack[8][0] ),
    .A2(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08790_ (.I(_02472_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08791_ (.A1(_02282_),
    .A2(_03034_),
    .B(_02489_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08792_ (.A1(_03001_),
    .A2(_03030_),
    .B1(_03033_),
    .B2(_03035_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08793_ (.I(_01830_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08794_ (.I(_01839_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08795_ (.A1(_03037_),
    .A2(_02488_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08796_ (.I(_03031_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08797_ (.I(_02481_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08798_ (.A1(\as2650.stack[8][1] ),
    .A2(_03039_),
    .B(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08799_ (.A1(_03036_),
    .A2(_03030_),
    .B1(_03038_),
    .B2(_03041_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(\as2650.stack[8][2] ),
    .A2(_03032_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08801_ (.A1(_03014_),
    .A2(_02483_),
    .B(_03040_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(_02441_),
    .A2(_03030_),
    .B1(_03042_),
    .B2(_03043_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_02298_),
    .A2(_03034_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08804_ (.A1(\as2650.stack[8][3] ),
    .A2(_03039_),
    .B(_03040_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08805_ (.A1(_02444_),
    .A2(_03030_),
    .B1(_03044_),
    .B2(_03045_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08806_ (.I(_02481_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08807_ (.A1(_02393_),
    .A2(_03034_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08808_ (.A1(\as2650.stack[8][4] ),
    .A2(_03039_),
    .B(_03040_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08809_ (.A1(_02688_),
    .A2(_03046_),
    .B1(_03047_),
    .B2(_03048_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08810_ (.A1(\as2650.stack[8][5] ),
    .A2(_03032_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08811_ (.A1(_03023_),
    .A2(_02483_),
    .B(_03029_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08812_ (.A1(_02453_),
    .A2(_03046_),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08813_ (.I(_01901_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(_02310_),
    .A2(_03034_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08815_ (.A1(\as2650.stack[8][6] ),
    .A2(_03039_),
    .B(_03029_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08816_ (.A1(_03051_),
    .A2(_03046_),
    .B1(_03052_),
    .B2(_03053_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(\as2650.stack[8][7] ),
    .A2(_03032_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08818_ (.A1(_02402_),
    .A2(_02483_),
    .B(_03029_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08819_ (.A1(_02459_),
    .A2(_03046_),
    .B1(_03054_),
    .B2(_03055_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08820_ (.I(_02344_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08821_ (.I(_03056_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08822_ (.A1(_02275_),
    .A2(_03004_),
    .A3(_02277_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08823_ (.I(_03058_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08824_ (.A1(\as2650.stack[11][0] ),
    .A2(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08825_ (.I(_01824_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08826_ (.I(_02338_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08827_ (.A1(_03061_),
    .A2(_03062_),
    .B(_02353_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08828_ (.A1(_03001_),
    .A2(_03057_),
    .B1(_03060_),
    .B2(_03063_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(_03037_),
    .A2(_02352_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08830_ (.I(_03058_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08831_ (.I(_02345_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08832_ (.A1(\as2650.stack[11][1] ),
    .A2(_03065_),
    .B(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08833_ (.A1(_03036_),
    .A2(_03057_),
    .B1(_03064_),
    .B2(_03067_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08834_ (.I(_01844_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(\as2650.stack[11][2] ),
    .A2(_03059_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08836_ (.A1(_03014_),
    .A2(_03062_),
    .B(_03066_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08837_ (.A1(_03068_),
    .A2(_03057_),
    .B1(_03069_),
    .B2(_03070_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08838_ (.I(_01862_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(\as2650.stack[11][3] ),
    .A2(_03059_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08840_ (.A1(_02388_),
    .A2(_02347_),
    .B(_03066_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08841_ (.A1(_03071_),
    .A2(_03057_),
    .B1(_03072_),
    .B2(_03073_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08842_ (.I(_02345_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08843_ (.I(_01883_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08844_ (.A1(_03075_),
    .A2(_03062_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08845_ (.A1(\as2650.stack[11][4] ),
    .A2(_03065_),
    .B(_03066_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08846_ (.A1(_02688_),
    .A2(_03074_),
    .B1(_03076_),
    .B2(_03077_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08847_ (.I(_01888_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08848_ (.A1(\as2650.stack[11][5] ),
    .A2(_03059_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08849_ (.A1(_03023_),
    .A2(_02347_),
    .B(_03056_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08850_ (.A1(_03078_),
    .A2(_03074_),
    .B1(_03079_),
    .B2(_03080_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(\as2650.stack[11][6] ),
    .A2(_03065_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08852_ (.A1(_02695_),
    .A2(_02347_),
    .B(_03056_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08853_ (.A1(_03051_),
    .A2(_03074_),
    .B1(_03081_),
    .B2(_03082_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08854_ (.I(_01913_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08855_ (.A1(_02314_),
    .A2(_03062_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08856_ (.A1(\as2650.stack[11][7] ),
    .A2(_03065_),
    .B(_03056_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08857_ (.A1(_03083_),
    .A2(_03074_),
    .B1(_03084_),
    .B2(_03085_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08858_ (.I(_02746_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08859_ (.I(_03086_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08860_ (.I(_02034_),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08861_ (.A1(_01798_),
    .A2(_03088_),
    .A3(_02427_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08862_ (.I(_03089_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08863_ (.A1(\as2650.stack[1][0] ),
    .A2(_03090_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08864_ (.A1(_02281_),
    .A2(_02749_),
    .B(_02747_),
    .C(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08865_ (.A1(_02372_),
    .A2(_03087_),
    .B(_03092_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08866_ (.I(_03089_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(\as2650.stack[1][1] ),
    .A2(_03093_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08868_ (.I(_02742_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08869_ (.A1(_02291_),
    .A2(_03095_),
    .B(_02755_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08870_ (.A1(_03036_),
    .A2(_03087_),
    .B1(_03094_),
    .B2(_03096_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08871_ (.A1(\as2650.stack[1][2] ),
    .A2(_03093_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08872_ (.I(_02747_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08873_ (.A1(_03014_),
    .A2(_03095_),
    .B(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08874_ (.A1(_03068_),
    .A2(_03087_),
    .B1(_03097_),
    .B2(_03099_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08875_ (.I(_01869_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08876_ (.A1(_03100_),
    .A2(_02754_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08877_ (.A1(\as2650.stack[1][3] ),
    .A2(_03090_),
    .B(_03098_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08878_ (.A1(_03071_),
    .A2(_03087_),
    .B1(_03101_),
    .B2(_03102_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08879_ (.I(_01459_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08880_ (.I(_03086_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(_03075_),
    .A2(_03095_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08882_ (.A1(\as2650.stack[1][4] ),
    .A2(_03090_),
    .B(_03098_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08883_ (.A1(_03103_),
    .A2(_03104_),
    .B1(_03105_),
    .B2(_03106_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08884_ (.A1(\as2650.stack[1][5] ),
    .A2(_03093_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08885_ (.A1(_03023_),
    .A2(_03095_),
    .B(_03098_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08886_ (.A1(_03078_),
    .A2(_03104_),
    .B1(_03107_),
    .B2(_03108_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08887_ (.A1(\as2650.stack[1][6] ),
    .A2(_03093_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08888_ (.A1(_02695_),
    .A2(_02749_),
    .B(_03086_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08889_ (.A1(_03051_),
    .A2(_03104_),
    .B1(_03109_),
    .B2(_03110_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08890_ (.A1(\as2650.stack[1][7] ),
    .A2(_03090_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08891_ (.I(_01921_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08892_ (.A1(_03112_),
    .A2(_02749_),
    .B(_03086_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08893_ (.A1(_03083_),
    .A2(_03104_),
    .B1(_03111_),
    .B2(_03113_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08894_ (.A1(_00995_),
    .A2(_00962_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08895_ (.I(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08896_ (.A1(_01027_),
    .A2(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08897_ (.A1(_00983_),
    .A2(_03115_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08898_ (.A1(_00968_),
    .A2(_00436_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08899_ (.A1(_01009_),
    .A2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08900_ (.A1(_01013_),
    .A2(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08901_ (.I(_03118_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08902_ (.A1(_01127_),
    .A2(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08903_ (.I(_03122_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08904_ (.A1(_00584_),
    .A2(_00991_),
    .A3(_00992_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08905_ (.A1(_01140_),
    .A2(_00972_),
    .A3(_03124_),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08906_ (.A1(_00999_),
    .A2(_03118_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08907_ (.I(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08908_ (.I(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08909_ (.A1(_03123_),
    .A2(_03125_),
    .A3(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08910_ (.A1(_03116_),
    .A2(_03117_),
    .A3(_03120_),
    .A4(_03129_),
    .Z(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08911_ (.I(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_00937_),
    .A2(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08913_ (.I(_03132_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08914_ (.I(_03117_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08915_ (.A1(_01140_),
    .A2(_00972_),
    .A3(_03124_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08916_ (.A1(_00536_),
    .A2(_00970_),
    .A3(_00974_),
    .A4(_00561_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08917_ (.A1(_01191_),
    .A2(_03136_),
    .A3(_03115_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08918_ (.A1(_01102_),
    .A2(_01104_),
    .A3(_03121_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08919_ (.I(_03138_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08920_ (.A1(_01113_),
    .A2(_03119_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08921_ (.I(_03140_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08922_ (.I(_03138_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08923_ (.A1(_01118_),
    .A2(_01119_),
    .A3(_03118_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08924_ (.I(_03140_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08925_ (.A1(_00449_),
    .A2(_03143_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08926_ (.A1(_02862_),
    .A2(_03143_),
    .B(_03144_),
    .C(_03145_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08927_ (.A1(_01111_),
    .A2(_03141_),
    .B(_03142_),
    .C(_03146_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08928_ (.A1(_01110_),
    .A2(_03139_),
    .B(_03147_),
    .C(_03123_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08929_ (.A1(_01006_),
    .A2(_03114_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08930_ (.I(_03149_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08931_ (.A1(_01100_),
    .A2(_03150_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08932_ (.A1(_03148_),
    .A2(_03151_),
    .B(_03137_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08933_ (.A1(_01098_),
    .A2(_03137_),
    .B(_03152_),
    .C(_03117_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08934_ (.A1(_01089_),
    .A2(_03134_),
    .B(_03135_),
    .C(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08935_ (.I(_03125_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(net80),
    .A2(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08937_ (.A1(_03154_),
    .A2(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(_01141_),
    .A2(_01126_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08939_ (.A1(_00926_),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08940_ (.A1(_00794_),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08941_ (.A1(_03160_),
    .A2(_03132_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08942_ (.I(_03161_),
    .Z(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08943_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_03162_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_03159_),
    .Z(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08945_ (.I(_03164_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08946_ (.A1(_01139_),
    .A2(_01151_),
    .A3(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08947_ (.A1(_03133_),
    .A2(_03157_),
    .B(_03163_),
    .C(_03166_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08948_ (.I(_03132_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08949_ (.I(_03125_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08950_ (.A1(_01191_),
    .A2(_03136_),
    .A3(_03115_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08951_ (.I(_03169_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08952_ (.A1(_01221_),
    .A2(_01222_),
    .A3(_03121_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08953_ (.I(_03126_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08954_ (.A1(_00451_),
    .A2(_03127_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08955_ (.A1(_01211_),
    .A2(_03172_),
    .B(_03144_),
    .C(_03173_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08956_ (.A1(_01204_),
    .A2(_03141_),
    .B(_03142_),
    .C(_03174_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08957_ (.A1(_01206_),
    .A2(_00637_),
    .A3(_03119_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08958_ (.I(_03149_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08959_ (.A1(_01217_),
    .A2(_03176_),
    .B(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08960_ (.A1(_01202_),
    .A2(_03150_),
    .B1(_03175_),
    .B2(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08961_ (.A1(_03169_),
    .A2(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08962_ (.A1(_01200_),
    .A2(_03170_),
    .B(_03171_),
    .C(_03180_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08963_ (.I(_03117_),
    .Z(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08964_ (.A1(_01229_),
    .A2(_03182_),
    .B(_03135_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08965_ (.A1(_03181_),
    .A2(_03183_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08966_ (.A1(_01188_),
    .A2(_03168_),
    .B(_03184_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08967_ (.A1(_01243_),
    .A2(_03165_),
    .B1(_03162_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03167_),
    .A2(_03185_),
    .B(_03186_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08969_ (.I(_00426_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08970_ (.I(_03144_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08971_ (.I(_03127_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08972_ (.I(_03140_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08973_ (.A1(_00443_),
    .A2(_03172_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08974_ (.A1(_02866_),
    .A2(_03189_),
    .B(_03190_),
    .C(_03191_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08975_ (.A1(_03187_),
    .A2(_03188_),
    .B(_03142_),
    .C(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08976_ (.A1(_01249_),
    .A2(_03176_),
    .B(_03177_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08977_ (.A1(_01246_),
    .A2(_03150_),
    .B1(_03193_),
    .B2(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08978_ (.A1(_03169_),
    .A2(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08979_ (.A1(_01269_),
    .A2(_03170_),
    .B(_03171_),
    .C(_03196_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08980_ (.A1(_01275_),
    .A2(_03182_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08981_ (.A1(_03197_),
    .A2(_03198_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08982_ (.A1(_01299_),
    .A2(_03155_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08983_ (.A1(_03168_),
    .A2(_03199_),
    .B(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08984_ (.I(_03164_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08985_ (.I(_03161_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08986_ (.A1(_01316_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(\as2650.r123_2[1][2] ),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08987_ (.A1(_03167_),
    .A2(_03201_),
    .B(_03204_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08988_ (.I(_03135_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08989_ (.I(_01367_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08990_ (.I(_03116_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08991_ (.I(_03207_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08992_ (.I(_03149_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08993_ (.I(_03176_),
    .Z(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08994_ (.A1(_00999_),
    .A2(_03121_),
    .B(_00428_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08995_ (.A1(_02871_),
    .A2(_03172_),
    .B(_03190_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08996_ (.A1(_01497_),
    .A2(_03141_),
    .B1(_03211_),
    .B2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08997_ (.A1(_03210_),
    .A2(_03213_),
    .B(_03123_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_01345_),
    .A2(_03210_),
    .B(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08999_ (.A1(_02132_),
    .A2(_03209_),
    .B(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(_03208_),
    .A2(_03216_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09001_ (.A1(_01362_),
    .A2(_03208_),
    .B(_03134_),
    .C(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09002_ (.A1(_03206_),
    .A2(_03134_),
    .B(_03205_),
    .C(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09003_ (.A1(_01343_),
    .A2(_03205_),
    .B(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09004_ (.A1(_01394_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(\as2650.r123_2[1][3] ),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09005_ (.A1(_03167_),
    .A2(_03220_),
    .B(_03221_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09006_ (.A1(_01428_),
    .A2(_03182_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09007_ (.A1(_01398_),
    .A2(_01401_),
    .A3(_01402_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09008_ (.A1(_00432_),
    .A2(_03128_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09009_ (.A1(_01409_),
    .A2(_03128_),
    .B(_03188_),
    .C(_03224_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09010_ (.A1(_01412_),
    .A2(_03188_),
    .B(_03139_),
    .C(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09011_ (.A1(_03187_),
    .A2(_03210_),
    .B(_03209_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09012_ (.A1(_01419_),
    .A2(_03209_),
    .B1(_03226_),
    .B2(_03227_),
    .C(_03207_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09013_ (.A1(_03223_),
    .A2(_03208_),
    .B(_03134_),
    .C(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09014_ (.A1(_03222_),
    .A2(_03229_),
    .B(_03155_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09015_ (.A1(_01456_),
    .A2(_03168_),
    .B(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09016_ (.I(_03231_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09017_ (.I(_01140_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09018_ (.A1(_03233_),
    .A2(_01460_),
    .A3(_01126_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09019_ (.A1(_01485_),
    .A2(_03234_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09020_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_03162_),
    .B(_03235_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09021_ (.A1(_03167_),
    .A2(_03232_),
    .B(_03236_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09022_ (.A1(_01496_),
    .A2(_03150_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09023_ (.A1(_02590_),
    .A2(_03189_),
    .B(_03190_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09024_ (.A1(_00425_),
    .A2(_03128_),
    .B(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09025_ (.A1(_01595_),
    .A2(_03188_),
    .B(_03139_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09026_ (.A1(_00429_),
    .A2(_03139_),
    .B1(_03239_),
    .B2(_03240_),
    .C(_03123_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09027_ (.A1(_03237_),
    .A2(_03241_),
    .B(_03207_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09028_ (.A1(_01509_),
    .A2(_03208_),
    .B(_03182_),
    .C(_03242_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09029_ (.I(_03171_),
    .Z(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09030_ (.A1(_01493_),
    .A2(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(_03243_),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09032_ (.A1(_01534_),
    .A2(_03155_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09033_ (.A1(_03168_),
    .A2(_03246_),
    .B(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09034_ (.A1(_01568_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(\as2650.r123_2[1][5] ),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09035_ (.A1(_03133_),
    .A2(_03248_),
    .B(_03249_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09036_ (.A1(_01575_),
    .A2(_03172_),
    .B(_03144_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09037_ (.A1(_00422_),
    .A2(_03189_),
    .B(_03250_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09038_ (.A1(_01109_),
    .A2(_03190_),
    .B(_03138_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09039_ (.A1(_01570_),
    .A2(_03142_),
    .B1(_03251_),
    .B2(_03252_),
    .C(_03122_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09040_ (.A1(_01583_),
    .A2(_03177_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09041_ (.A1(_03253_),
    .A2(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09042_ (.A1(_03169_),
    .A2(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09043_ (.A1(_01592_),
    .A2(_03170_),
    .B(_03171_),
    .C(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09044_ (.A1(_01597_),
    .A2(_03244_),
    .B(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09045_ (.I0(_01622_),
    .I1(_03258_),
    .S(_03205_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_01667_),
    .A2(_03234_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09047_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_03162_),
    .B(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09048_ (.A1(_03133_),
    .A2(_03259_),
    .B(_03261_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09049_ (.A1(_00832_),
    .A2(_03127_),
    .B(_03140_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09050_ (.A1(_05840_),
    .A2(_03189_),
    .B(_03262_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09051_ (.A1(_01673_),
    .A2(_03141_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09052_ (.A1(_03176_),
    .A2(_03263_),
    .A3(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09053_ (.A1(_02886_),
    .A2(_03210_),
    .B(_03265_),
    .C(_03177_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09054_ (.A1(_01916_),
    .A2(_03209_),
    .B(_03266_),
    .C(_03207_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09055_ (.A1(_01687_),
    .A2(_03170_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09056_ (.A1(_03267_),
    .A2(_03268_),
    .B(_03244_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09057_ (.A1(_01692_),
    .A2(_03244_),
    .B(_03269_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09058_ (.I0(_01717_),
    .I1(_03270_),
    .S(_03135_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09059_ (.A1(_01758_),
    .A2(_03202_),
    .B1(_03203_),
    .B2(\as2650.r123_2[1][7] ),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09060_ (.A1(_03133_),
    .A2(_03271_),
    .B(_03272_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09061_ (.I(\as2650.r123_2[0][0] ),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09062_ (.A1(_00936_),
    .A2(_01928_),
    .B(_03158_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09063_ (.A1(_00955_),
    .A2(_03130_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09064_ (.A1(_00513_),
    .A2(_03274_),
    .A3(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09065_ (.I(_03276_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09066_ (.I(_03277_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09067_ (.I(_03157_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09068_ (.I(_03275_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09069_ (.A1(_01940_),
    .A2(_03158_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09070_ (.I(_03281_),
    .Z(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09071_ (.I(_03282_),
    .Z(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09072_ (.A1(_03159_),
    .A2(_03274_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09073_ (.I(_03284_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09074_ (.I(_03281_),
    .Z(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09075_ (.A1(_01137_),
    .A2(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09076_ (.A1(_02011_),
    .A2(_03283_),
    .B(_03285_),
    .C(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09077_ (.A1(_03279_),
    .A2(_03280_),
    .B(_03277_),
    .C(_03288_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09078_ (.A1(_03273_),
    .A2(_03278_),
    .B(_03289_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09079_ (.I(\as2650.r123_2[0][1] ),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09080_ (.I(_03185_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09081_ (.I(_03276_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09082_ (.A1(_01240_),
    .A2(_03286_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09083_ (.A1(_02056_),
    .A2(_03283_),
    .B(_03285_),
    .C(_03293_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09084_ (.A1(_03291_),
    .A2(_03280_),
    .B(_03292_),
    .C(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09085_ (.A1(_03290_),
    .A2(_03278_),
    .B(_03295_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09086_ (.I(\as2650.r123_2[0][2] ),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09087_ (.I(_03201_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09088_ (.I(_03281_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09089_ (.I(_03284_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09090_ (.A1(_01247_),
    .A2(_03286_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09091_ (.A1(_02096_),
    .A2(_03298_),
    .B(_03299_),
    .C(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09092_ (.A1(_03297_),
    .A2(_03280_),
    .B(_03292_),
    .C(_03301_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09093_ (.A1(_03296_),
    .A2(_03278_),
    .B(_03302_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09094_ (.I(\as2650.r123_2[0][3] ),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09095_ (.I(_03277_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09096_ (.A1(_02133_),
    .A2(_03286_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09097_ (.A1(_02131_),
    .A2(_03283_),
    .B(_03285_),
    .C(_03305_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09098_ (.A1(_03277_),
    .A2(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09099_ (.A1(_01343_),
    .A2(_03205_),
    .B(_03219_),
    .C(_03280_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09100_ (.A1(_03303_),
    .A2(_03304_),
    .B1(_03307_),
    .B2(_03308_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09101_ (.I(\as2650.r123_2[0][4] ),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09102_ (.I(_03275_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09103_ (.A1(_02156_),
    .A2(_03282_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09104_ (.A1(_02155_),
    .A2(_03298_),
    .B(_03299_),
    .C(_03311_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09105_ (.A1(_03231_),
    .A2(_03310_),
    .B(_03292_),
    .C(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09106_ (.A1(_03309_),
    .A2(_03278_),
    .B(_03313_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09107_ (.I(\as2650.r123_2[0][5] ),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09108_ (.I(_03248_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09109_ (.I(_01896_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09110_ (.A1(_03316_),
    .A2(_03282_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09111_ (.A1(_02176_),
    .A2(_03298_),
    .B(_03299_),
    .C(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09112_ (.A1(_03315_),
    .A2(_03310_),
    .B(_03292_),
    .C(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09113_ (.A1(_03314_),
    .A2(_03304_),
    .B(_03319_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09114_ (.I(\as2650.r123_2[0][6] ),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09115_ (.I(_03259_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09116_ (.A1(_01908_),
    .A2(_03282_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09117_ (.A1(_02193_),
    .A2(_03298_),
    .B(_03299_),
    .C(_03322_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09118_ (.A1(_03321_),
    .A2(_03310_),
    .B(_03276_),
    .C(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09119_ (.A1(_03320_),
    .A2(_03304_),
    .B(_03324_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09120_ (.I(\as2650.r123_2[0][7] ),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09121_ (.I(_03271_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09122_ (.A1(_02199_),
    .A2(_03283_),
    .A3(_03285_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09123_ (.A1(_03326_),
    .A2(_03310_),
    .B(_03276_),
    .C(_03327_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09124_ (.A1(_03325_),
    .A2(_03304_),
    .B(_03328_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09125_ (.I(_02498_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09126_ (.I(_03329_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09127_ (.I(_02112_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09128_ (.A1(_02703_),
    .A2(_01781_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09129_ (.A1(_02666_),
    .A2(_03331_),
    .A3(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09130_ (.I(_03333_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09131_ (.A1(\as2650.stack[7][0] ),
    .A2(_03334_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09132_ (.I(_02494_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09133_ (.A1(_03061_),
    .A2(_03336_),
    .B(_02507_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09134_ (.A1(_03001_),
    .A2(_03330_),
    .B1(_03335_),
    .B2(_03337_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09135_ (.I(_03333_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09136_ (.A1(\as2650.stack[7][1] ),
    .A2(_03338_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09137_ (.A1(_02380_),
    .A2(_02501_),
    .B(_02499_),
    .C(_03339_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09138_ (.A1(_01832_),
    .A2(_03330_),
    .B(_03340_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09139_ (.A1(\as2650.stack[7][2] ),
    .A2(_03334_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09140_ (.I(_01857_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09141_ (.I(_02499_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09142_ (.A1(_03342_),
    .A2(_03336_),
    .B(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09143_ (.A1(_03068_),
    .A2(_03330_),
    .B1(_03341_),
    .B2(_03344_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09144_ (.A1(_03100_),
    .A2(_02506_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09145_ (.A1(\as2650.stack[7][3] ),
    .A2(_03338_),
    .B(_03343_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09146_ (.A1(_03071_),
    .A2(_03330_),
    .B1(_03345_),
    .B2(_03346_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09147_ (.I(_03329_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09148_ (.A1(_03075_),
    .A2(_03336_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09149_ (.A1(\as2650.stack[7][4] ),
    .A2(_03338_),
    .B(_03343_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09150_ (.A1(_03103_),
    .A2(_03347_),
    .B1(_03348_),
    .B2(_03349_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09151_ (.A1(\as2650.stack[7][5] ),
    .A2(_03334_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09152_ (.I(_01898_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09153_ (.A1(_03351_),
    .A2(_03336_),
    .B(_03343_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09154_ (.A1(_03078_),
    .A2(_03347_),
    .B1(_03350_),
    .B2(_03352_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(\as2650.stack[7][6] ),
    .A2(_03334_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09156_ (.I(_01910_),
    .Z(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09157_ (.A1(_03354_),
    .A2(_02501_),
    .B(_03329_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09158_ (.A1(_03051_),
    .A2(_03347_),
    .B1(_03353_),
    .B2(_03355_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(\as2650.stack[7][7] ),
    .A2(_03338_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09160_ (.A1(_03112_),
    .A2(_02501_),
    .B(_03329_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09161_ (.A1(_03083_),
    .A2(_03347_),
    .B1(_03356_),
    .B2(_03357_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09162_ (.A1(_00479_),
    .A2(_03131_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09163_ (.I(_03358_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09164_ (.I(_03359_),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09165_ (.A1(_03160_),
    .A2(_03358_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09166_ (.I(_03361_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09168_ (.I(_03164_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09169_ (.A1(_01726_),
    .A2(_01756_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09170_ (.A1(_01726_),
    .A2(_01756_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09171_ (.A1(_01721_),
    .A2(_03365_),
    .B(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09172_ (.A1(_01738_),
    .A2(_01754_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09173_ (.A1(_01732_),
    .A2(_03368_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09174_ (.A1(_01729_),
    .A2(_01755_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09175_ (.A1(_03369_),
    .A2(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09176_ (.A1(_01323_),
    .A2(_01634_),
    .A3(_01736_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09177_ (.A1(_01734_),
    .A2(_01735_),
    .B(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09178_ (.A1(_01740_),
    .A2(_01753_),
    .Z(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09179_ (.A1(_01738_),
    .A2(_01754_),
    .B(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09180_ (.A1(_05817_),
    .A2(_01653_),
    .A3(_01654_),
    .A4(_01751_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09181_ (.A1(_01745_),
    .A2(_01752_),
    .B(_03376_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09182_ (.A1(_05737_),
    .A2(_01647_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09183_ (.A1(_05737_),
    .A2(_01235_),
    .B1(_02254_),
    .B2(_01305_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09184_ (.A1(_01306_),
    .A2(_03378_),
    .B(_03379_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09185_ (.A1(_01660_),
    .A2(_01749_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09186_ (.A1(_01747_),
    .A2(_01750_),
    .B(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(\as2650.r0[1] ),
    .A2(_01748_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09188_ (.A1(\as2650.r0[5] ),
    .A2(_01380_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(_05830_),
    .A2(_01310_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09190_ (.A1(_03383_),
    .A2(_03384_),
    .A3(_03385_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09191_ (.A1(_03382_),
    .A2(_03386_),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09192_ (.A1(_03380_),
    .A2(_03387_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09193_ (.A1(_03377_),
    .A2(_03388_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09194_ (.A1(_01742_),
    .A2(_01743_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09195_ (.A1(_01741_),
    .A2(_01744_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09196_ (.A1(_03390_),
    .A2(_03391_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(_05778_),
    .A2(_01629_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09198_ (.A1(_03392_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09199_ (.A1(_01417_),
    .A2(_01467_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09200_ (.A1(_03394_),
    .A2(_03395_),
    .Z(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09201_ (.A1(_03389_),
    .A2(_03396_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09202_ (.A1(_03375_),
    .A2(_03397_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09203_ (.A1(_03373_),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09204_ (.A1(_03371_),
    .A2(_03399_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09205_ (.A1(_03367_),
    .A2(_03400_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09206_ (.A1(_03364_),
    .A2(_03401_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09207_ (.A1(_03157_),
    .A2(_03360_),
    .B(_03363_),
    .C(_03402_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09208_ (.A1(_03371_),
    .A2(_03399_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09209_ (.A1(_03367_),
    .A2(_03400_),
    .B(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(_03375_),
    .A2(_03397_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09211_ (.A1(_03373_),
    .A2(_03398_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09212_ (.A1(_03405_),
    .A2(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09213_ (.A1(_03392_),
    .A2(_03393_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09214_ (.A1(_03394_),
    .A2(_03395_),
    .B(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_03377_),
    .A2(_03388_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_03389_),
    .A2(_03396_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(_03410_),
    .A2(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(_03380_),
    .A2(_03387_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09219_ (.A1(_03382_),
    .A2(_03386_),
    .B(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_01374_),
    .A2(_02254_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09221_ (.I(_01748_),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(_05758_),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09223_ (.A1(_03383_),
    .A2(_03384_),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09224_ (.A1(_01479_),
    .A2(_03417_),
    .B1(_03418_),
    .B2(_03385_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(\as2650.r0[2] ),
    .A2(_01748_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09226_ (.A1(\as2650.r0[6] ),
    .A2(_01379_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09227_ (.A1(_03420_),
    .A2(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09228_ (.A1(\as2650.r0[7] ),
    .A2(_01310_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09229_ (.A1(_03422_),
    .A2(_03423_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09230_ (.A1(_03419_),
    .A2(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09231_ (.A1(_03415_),
    .A2(_03425_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09232_ (.I(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09233_ (.A1(_03414_),
    .A2(_03427_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_01306_),
    .A2(_03378_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_05769_),
    .A2(_01629_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09236_ (.A1(_05760_),
    .A2(_01467_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09237_ (.A1(_03429_),
    .A2(_03430_),
    .A3(_03431_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09238_ (.I(_03432_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09239_ (.A1(_03428_),
    .A2(_03433_),
    .Z(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09240_ (.A1(_03412_),
    .A2(_03434_),
    .Z(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09241_ (.A1(_03409_),
    .A2(_03435_),
    .Z(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09242_ (.A1(_03407_),
    .A2(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09243_ (.A1(_03404_),
    .A2(_03437_),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(_03364_),
    .A2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09245_ (.I(_03361_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09246_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09247_ (.A1(_03185_),
    .A2(_03360_),
    .B(_03439_),
    .C(_03441_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(_03407_),
    .A2(_03436_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09249_ (.A1(_03404_),
    .A2(_03437_),
    .B(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09250_ (.A1(_03412_),
    .A2(_03434_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09251_ (.A1(_03409_),
    .A2(_03435_),
    .B(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09252_ (.A1(_03429_),
    .A2(_03430_),
    .Z(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09253_ (.A1(_03429_),
    .A2(_03430_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09254_ (.A1(_03446_),
    .A2(_03431_),
    .B(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09255_ (.A1(_03414_),
    .A2(_03427_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(_03428_),
    .A2(_03433_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09257_ (.A1(_03449_),
    .A2(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(_05832_),
    .A2(_01633_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09259_ (.A1(_01495_),
    .A2(_01630_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_05832_),
    .A2(_01630_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09261_ (.A1(_03431_),
    .A2(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09262_ (.A1(_03452_),
    .A2(_03453_),
    .B(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_03419_),
    .A2(_03424_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09264_ (.A1(_01323_),
    .A2(_02255_),
    .A3(_03425_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(_03457_),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09266_ (.A1(_05737_),
    .A2(_03416_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09267_ (.A1(_01656_),
    .A2(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09268_ (.I(_03416_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09269_ (.A1(_05738_),
    .A2(_01381_),
    .B1(_03462_),
    .B2(_01373_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09270_ (.A1(_03461_),
    .A2(_03463_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09271_ (.A1(_05831_),
    .A2(_03416_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09272_ (.A1(_01554_),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09273_ (.A1(_03422_),
    .A2(_03423_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09274_ (.A1(_03466_),
    .A2(_03467_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09275_ (.A1(_03464_),
    .A2(_03468_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(_01417_),
    .A2(_02254_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09277_ (.A1(_03469_),
    .A2(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09278_ (.A1(_03459_),
    .A2(_03471_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09279_ (.A1(_03456_),
    .A2(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09280_ (.A1(_03451_),
    .A2(_03473_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09281_ (.A1(_03448_),
    .A2(_03474_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09282_ (.A1(_03445_),
    .A2(_03475_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09283_ (.A1(_03443_),
    .A2(_03476_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(_03364_),
    .A2(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_03440_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09286_ (.A1(_03201_),
    .A2(_03360_),
    .B(_03478_),
    .C(_03479_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09287_ (.A1(_03445_),
    .A2(_03475_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09288_ (.A1(_03443_),
    .A2(_03476_),
    .B(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(_03451_),
    .A2(_03473_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09290_ (.A1(_03448_),
    .A2(_03474_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(_03459_),
    .A2(_03471_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09292_ (.A1(_03456_),
    .A2(_03472_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(_03484_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(_01676_),
    .A2(_01633_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09295_ (.A1(_05738_),
    .A2(_01630_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09296_ (.A1(_03452_),
    .A2(_03488_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09297_ (.I(_03489_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09298_ (.A1(_03454_),
    .A2(_03487_),
    .B(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09299_ (.A1(_01418_),
    .A2(_02256_),
    .A3(_03469_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09300_ (.A1(_03464_),
    .A2(_03468_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09301_ (.A1(_05769_),
    .A2(_03462_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(_01417_),
    .A2(_03461_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09303_ (.A1(_03494_),
    .A2(_03461_),
    .B(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09304_ (.A1(_05760_),
    .A2(_02255_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09305_ (.A1(_03496_),
    .A2(_03497_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09306_ (.A1(_03493_),
    .A2(_03498_),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09307_ (.A1(_03491_),
    .A2(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09308_ (.A1(_03486_),
    .A2(_03500_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09309_ (.A1(_03455_),
    .A2(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09310_ (.A1(_03482_),
    .A2(_03483_),
    .B(_03502_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09311_ (.A1(_03482_),
    .A2(_03483_),
    .A3(_03502_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09312_ (.A1(_03503_),
    .A2(_03504_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09313_ (.A1(_03481_),
    .A2(_03505_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09314_ (.A1(_03364_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_03440_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09316_ (.A1(_03220_),
    .A2(_03360_),
    .B(_03507_),
    .C(_03508_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09317_ (.A1(_03486_),
    .A2(_03500_),
    .B1(_03501_),
    .B2(_03455_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09318_ (.A1(_03493_),
    .A2(_03498_),
    .B1(_03499_),
    .B2(_03491_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09319_ (.A1(_05831_),
    .A2(_02255_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09320_ (.A1(_03417_),
    .A2(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09321_ (.A1(_03496_),
    .A2(_03497_),
    .B(_03495_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09322_ (.A1(_03512_),
    .A2(_03513_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09323_ (.A1(_03488_),
    .A2(_03514_),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09324_ (.A1(_03510_),
    .A2(_03515_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09325_ (.A1(_03489_),
    .A2(_03516_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09326_ (.A1(_03509_),
    .A2(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09327_ (.A1(_03443_),
    .A2(_03476_),
    .B(_03503_),
    .C(_03480_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09328_ (.A1(_03504_),
    .A2(_03519_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09329_ (.A1(_03518_),
    .A2(_03520_),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09330_ (.I(_03358_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09331_ (.A1(_03231_),
    .A2(_03522_),
    .B1(_03362_),
    .B2(\as2650.r123_2[2][4] ),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09332_ (.A1(_03234_),
    .A2(_03521_),
    .B(_03523_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09333_ (.A1(_03504_),
    .A2(_03518_),
    .A3(_03519_),
    .B1(_03509_),
    .B2(_03517_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(_03512_),
    .A2(_03513_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09335_ (.A1(_01677_),
    .A2(_01631_),
    .A3(_03514_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09336_ (.A1(_03525_),
    .A2(_03526_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(_01676_),
    .A2(_02256_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09338_ (.A1(_01582_),
    .A2(_03462_),
    .A3(_03497_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09339_ (.A1(_03528_),
    .A2(_03529_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09340_ (.A1(_03527_),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09341_ (.A1(_03510_),
    .A2(_03515_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09342_ (.A1(_03490_),
    .A2(_03516_),
    .B(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09343_ (.A1(_03524_),
    .A2(_03531_),
    .A3(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(_03165_),
    .A2(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09345_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_03440_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09346_ (.A1(_03248_),
    .A2(_03359_),
    .B(_03535_),
    .C(_03536_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09347_ (.A1(_03531_),
    .A2(_03533_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09348_ (.A1(_03531_),
    .A2(_03533_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09349_ (.A1(_03524_),
    .A2(_03537_),
    .B(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(_03527_),
    .A2(_03530_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09351_ (.A1(_01916_),
    .A2(_03465_),
    .A3(_03497_),
    .B1(_03511_),
    .B2(_03460_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09352_ (.A1(_03540_),
    .A2(_03541_),
    .Z(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09353_ (.A1(_03539_),
    .A2(_03542_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09354_ (.A1(_03165_),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09355_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_03362_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09356_ (.A1(_03259_),
    .A2(_03359_),
    .B(_03544_),
    .C(_03545_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09357_ (.A1(_03528_),
    .A2(_03465_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09358_ (.A1(_03460_),
    .A2(_03511_),
    .A3(_03540_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09359_ (.A1(_03539_),
    .A2(_03542_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09360_ (.A1(_03546_),
    .A2(_03547_),
    .A3(_03548_),
    .B(_03164_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09361_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_03362_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09362_ (.A1(_03271_),
    .A2(_03359_),
    .B(_03549_),
    .C(_03550_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09363_ (.I(_02705_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09364_ (.I(_03551_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09365_ (.A1(_02666_),
    .A2(_03331_),
    .A3(_02427_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09366_ (.I(_03553_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09367_ (.A1(\as2650.stack[3][0] ),
    .A2(_03554_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09368_ (.A1(_02281_),
    .A2(_02708_),
    .B(_03551_),
    .C(_03555_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09369_ (.A1(_02372_),
    .A2(_03552_),
    .B(_03556_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09370_ (.I(_03553_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09371_ (.A1(\as2650.stack[3][1] ),
    .A2(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09372_ (.A1(_02380_),
    .A2(_02713_),
    .B(_02714_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09373_ (.A1(_03036_),
    .A2(_03552_),
    .B1(_03558_),
    .B2(_03559_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09374_ (.A1(\as2650.stack[3][2] ),
    .A2(_03557_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09375_ (.I(_02699_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09376_ (.I(_02706_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09377_ (.A1(_03342_),
    .A2(_03561_),
    .B(_03562_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09378_ (.A1(_03068_),
    .A2(_03552_),
    .B1(_03560_),
    .B2(_03563_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09379_ (.I(_03551_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09380_ (.A1(\as2650.stack[3][3] ),
    .A2(_03557_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09381_ (.A1(_02388_),
    .A2(_03561_),
    .B(_03562_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09382_ (.A1(_03071_),
    .A2(_03564_),
    .B1(_03565_),
    .B2(_03566_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09383_ (.A1(\as2650.stack[3][4] ),
    .A2(_03557_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09384_ (.A1(_02392_),
    .A2(_03561_),
    .B(_03562_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09385_ (.A1(_03103_),
    .A2(_03564_),
    .B1(_03567_),
    .B2(_03568_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09386_ (.A1(\as2650.stack[3][5] ),
    .A2(_03554_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09387_ (.A1(_03351_),
    .A2(_03561_),
    .B(_03562_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09388_ (.A1(_03078_),
    .A2(_03564_),
    .B1(_03569_),
    .B2(_03570_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09389_ (.A1(\as2650.stack[3][6] ),
    .A2(_03554_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09390_ (.A1(_01911_),
    .A2(_02708_),
    .B(_02706_),
    .C(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09391_ (.A1(_01903_),
    .A2(_03552_),
    .B(_03572_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09392_ (.A1(\as2650.stack[3][7] ),
    .A2(_03554_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09393_ (.A1(_03112_),
    .A2(_02708_),
    .B(_03551_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09394_ (.A1(_03083_),
    .A2(_03564_),
    .B1(_03573_),
    .B2(_03574_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09395_ (.I(_01760_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09396_ (.I(_02633_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09397_ (.I(_03576_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09398_ (.A1(_02666_),
    .A2(_03088_),
    .A3(_03332_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09399_ (.I(_03578_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09400_ (.A1(\as2650.stack[5][0] ),
    .A2(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09401_ (.A1(_03061_),
    .A2(_02641_),
    .B(_02642_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09402_ (.A1(_03575_),
    .A2(_03577_),
    .B1(_03580_),
    .B2(_03581_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09403_ (.I(_03578_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09404_ (.A1(\as2650.stack[5][1] ),
    .A2(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09405_ (.A1(_01839_),
    .A2(_02636_),
    .B(_02634_),
    .C(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09406_ (.A1(_02289_),
    .A2(_03577_),
    .B(_03584_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(\as2650.stack[5][2] ),
    .A2(_03579_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09408_ (.I(_02629_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09409_ (.I(_02634_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09410_ (.A1(_03342_),
    .A2(_03586_),
    .B(_03587_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09411_ (.A1(_01845_),
    .A2(_03577_),
    .B1(_03585_),
    .B2(_03588_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09412_ (.I(_01861_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(\as2650.stack[5][3] ),
    .A2(_03579_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09414_ (.A1(_01870_),
    .A2(_03586_),
    .B(_03587_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09415_ (.A1(_03589_),
    .A2(_03577_),
    .B1(_03590_),
    .B2(_03591_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09416_ (.I(_03576_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(\as2650.stack[5][4] ),
    .A2(_03579_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09418_ (.A1(_02392_),
    .A2(_03586_),
    .B(_03587_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09419_ (.A1(_03103_),
    .A2(_03592_),
    .B1(_03593_),
    .B2(_03594_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09420_ (.A1(\as2650.stack[5][5] ),
    .A2(_03582_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09421_ (.A1(_03351_),
    .A2(_03586_),
    .B(_03587_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09422_ (.A1(_01889_),
    .A2(_03592_),
    .B1(_03595_),
    .B2(_03596_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(\as2650.stack[5][6] ),
    .A2(_03582_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09424_ (.A1(_03354_),
    .A2(_02636_),
    .B(_03576_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09425_ (.A1(_01902_),
    .A2(_03592_),
    .B1(_03597_),
    .B2(_03598_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09426_ (.I(_01913_),
    .Z(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09427_ (.A1(\as2650.stack[5][7] ),
    .A2(_03582_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09428_ (.A1(_03112_),
    .A2(_02636_),
    .B(_03576_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09429_ (.A1(_03599_),
    .A2(_03592_),
    .B1(_03600_),
    .B2(_03601_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09430_ (.I(_02651_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09431_ (.I(_03602_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09432_ (.A1(_02424_),
    .A2(_02425_),
    .A3(_03332_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09433_ (.I(_03604_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09434_ (.A1(\as2650.stack[4][0] ),
    .A2(_03605_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09435_ (.I(_02646_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09436_ (.I(_02652_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09437_ (.A1(_03061_),
    .A2(_03607_),
    .B(_03608_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09438_ (.A1(_03575_),
    .A2(_03603_),
    .B1(_03606_),
    .B2(_03609_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09439_ (.A1(_03037_),
    .A2(_02659_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09440_ (.A1(\as2650.stack[4][1] ),
    .A2(_03605_),
    .B(_03608_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09441_ (.A1(_01831_),
    .A2(_03603_),
    .B1(_03610_),
    .B2(_03611_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09442_ (.I(_02652_),
    .Z(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09443_ (.A1(\as2650.stack[4][2] ),
    .A2(_02661_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09444_ (.I(_03604_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09445_ (.A1(_01858_),
    .A2(_03614_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(net49),
    .A2(_03612_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09447_ (.A1(_03612_),
    .A2(_03613_),
    .A3(_03615_),
    .B(_03616_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(\as2650.stack[4][3] ),
    .A2(_03605_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09449_ (.A1(_01870_),
    .A2(_03607_),
    .B(_03602_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09450_ (.A1(_03589_),
    .A2(_03603_),
    .B1(_03617_),
    .B2(_03618_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(_03075_),
    .A2(_03607_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09452_ (.A1(\as2650.stack[4][4] ),
    .A2(_03614_),
    .B(_03602_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09453_ (.A1(_01873_),
    .A2(_03603_),
    .B1(_03619_),
    .B2(_03620_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09454_ (.A1(\as2650.stack[4][5] ),
    .A2(_02661_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09455_ (.A1(_01899_),
    .A2(_03614_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09456_ (.A1(net52),
    .A2(_03608_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09457_ (.A1(_03612_),
    .A2(_03621_),
    .A3(_03622_),
    .B(_03623_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09458_ (.A1(\as2650.stack[4][6] ),
    .A2(_02647_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09459_ (.A1(_01911_),
    .A2(_03614_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(_02897_),
    .A2(_03608_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09461_ (.A1(_03612_),
    .A2(_03624_),
    .A3(_03625_),
    .B(_03626_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(\as2650.stack[4][7] ),
    .A2(_03605_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09463_ (.A1(_01922_),
    .A2(_03607_),
    .B(_03602_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09464_ (.A1(_03599_),
    .A2(_02653_),
    .B1(_03627_),
    .B2(_03628_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09465_ (.I(_02626_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09466_ (.I(_02603_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09467_ (.I(_02608_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09468_ (.I(\as2650.stack[6][0] ),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09469_ (.A1(_03632_),
    .A2(_02620_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09470_ (.A1(_02281_),
    .A2(_03630_),
    .B(_03631_),
    .C(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09471_ (.A1(_01761_),
    .A2(_03629_),
    .B(_03634_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09472_ (.A1(net86),
    .A2(_02626_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09473_ (.I(_02608_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09474_ (.A1(_02678_),
    .A2(_02604_),
    .B(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09475_ (.A1(\as2650.stack[6][1] ),
    .A2(_02621_),
    .B(_03637_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09476_ (.A1(_03635_),
    .A2(_03638_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09477_ (.I(\as2650.stack[6][2] ),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09478_ (.A1(_03639_),
    .A2(_02620_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09479_ (.A1(_01858_),
    .A2(_03630_),
    .B(_03631_),
    .C(_03640_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09480_ (.A1(_01846_),
    .A2(_03629_),
    .B(_03641_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09481_ (.I(\as2650.stack[6][3] ),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09482_ (.I(_02602_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09483_ (.A1(_03642_),
    .A2(_03643_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09484_ (.A1(_01870_),
    .A2(_03630_),
    .B(_03631_),
    .C(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09485_ (.A1(_01863_),
    .A2(_03629_),
    .B(_03645_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09486_ (.A1(_03233_),
    .A2(_02626_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09487_ (.I(_02156_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(_01880_),
    .A2(_02669_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09489_ (.A1(_03647_),
    .A2(_02669_),
    .B(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09490_ (.A1(_03649_),
    .A2(_02620_),
    .B(_03636_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(\as2650.stack[6][4] ),
    .A2(_03630_),
    .B(_03650_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(_03646_),
    .A2(_03651_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09493_ (.I(\as2650.stack[6][5] ),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09494_ (.A1(_03652_),
    .A2(_03643_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09495_ (.A1(_01899_),
    .A2(_02611_),
    .B(_03631_),
    .C(_03653_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09496_ (.A1(_01890_),
    .A2(_03629_),
    .B(_03654_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09497_ (.I(\as2650.stack[6][6] ),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09498_ (.A1(_03655_),
    .A2(_03643_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09499_ (.A1(_01911_),
    .A2(_02611_),
    .B(_03636_),
    .C(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09500_ (.A1(_01903_),
    .A2(_02609_),
    .B(_03657_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09501_ (.I(\as2650.stack[6][7] ),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09502_ (.A1(_03658_),
    .A2(_03643_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09503_ (.A1(_01922_),
    .A2(_02611_),
    .B(_03636_),
    .C(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09504_ (.A1(_01914_),
    .A2(_02609_),
    .B(_03660_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09505_ (.A1(_00797_),
    .A2(_02559_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09506_ (.A1(_00794_),
    .A2(_00917_),
    .A3(_02532_),
    .A4(_03661_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09507_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09508_ (.I0(\as2650.ivec[0] ),
    .I1(_01139_),
    .S(_03663_),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09509_ (.I(_03664_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09510_ (.I0(\as2650.ivec[1] ),
    .I1(_02676_),
    .S(_03663_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09511_ (.I(_03665_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09512_ (.I(_03662_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09513_ (.I(_03666_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09514_ (.A1(\as2650.ivec[2] ),
    .A2(_03667_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09515_ (.A1(_01847_),
    .A2(_03667_),
    .B(_03668_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09516_ (.A1(\as2650.ivec[3] ),
    .A2(_03663_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09517_ (.A1(_01354_),
    .A2(_03667_),
    .B(_03669_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09518_ (.I0(\as2650.ivec[4] ),
    .I1(_03647_),
    .S(_03666_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09519_ (.I(_03670_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09520_ (.I0(\as2650.ivec[5] ),
    .I1(_03316_),
    .S(_03666_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09521_ (.I(_03671_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09522_ (.I(_01908_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09523_ (.I0(\as2650.ivec[6] ),
    .I1(_03672_),
    .S(_03666_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09524_ (.I(_03673_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09525_ (.A1(\as2650.ivec[7] ),
    .A2(_03663_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09526_ (.A1(_02199_),
    .A2(_03667_),
    .B(_03674_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09527_ (.I(_02723_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09528_ (.I(_03675_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09529_ (.A1(_02275_),
    .A2(_02276_),
    .A3(_02427_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09530_ (.I(_03677_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09531_ (.A1(\as2650.stack[2][0] ),
    .A2(_03678_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09532_ (.I(_02719_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09533_ (.A1(_01825_),
    .A2(_03680_),
    .B(_02736_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09534_ (.A1(_03575_),
    .A2(_03676_),
    .B1(_03679_),
    .B2(_03681_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(\as2650.stack[2][1] ),
    .A2(_03678_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09536_ (.I(_02724_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09537_ (.A1(_02380_),
    .A2(_03680_),
    .B(_03683_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09538_ (.A1(_01831_),
    .A2(_03676_),
    .B1(_03682_),
    .B2(_03684_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09539_ (.A1(\as2650.stack[2][2] ),
    .A2(_03678_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09540_ (.A1(_03342_),
    .A2(_03680_),
    .B(_03683_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09541_ (.A1(_01845_),
    .A2(_03676_),
    .B1(_03685_),
    .B2(_03686_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(_03100_),
    .A2(_02735_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09543_ (.I(_03677_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09544_ (.A1(\as2650.stack[2][3] ),
    .A2(_03688_),
    .B(_03683_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09545_ (.A1(_03589_),
    .A2(_03676_),
    .B1(_03687_),
    .B2(_03689_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09546_ (.I(_02724_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09547_ (.A1(_01884_),
    .A2(_03680_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09548_ (.A1(\as2650.stack[2][4] ),
    .A2(_03688_),
    .B(_03683_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09549_ (.A1(_01873_),
    .A2(_03690_),
    .B1(_03691_),
    .B2(_03692_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(\as2650.stack[2][5] ),
    .A2(_03678_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09551_ (.A1(_03351_),
    .A2(_02727_),
    .B(_03675_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09552_ (.A1(_01889_),
    .A2(_03690_),
    .B1(_03693_),
    .B2(_03694_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09553_ (.A1(\as2650.stack[2][6] ),
    .A2(_03688_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09554_ (.A1(_03354_),
    .A2(_02727_),
    .B(_03675_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09555_ (.A1(_01902_),
    .A2(_03690_),
    .B1(_03695_),
    .B2(_03696_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(\as2650.stack[2][7] ),
    .A2(_03688_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09557_ (.A1(_01922_),
    .A2(_02727_),
    .B(_03675_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09558_ (.A1(_03599_),
    .A2(_03690_),
    .B1(_03697_),
    .B2(_03698_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(_00886_),
    .A2(_00878_),
    .B(_02859_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09560_ (.A1(_00462_),
    .A2(_00893_),
    .A3(_02783_),
    .A4(_02785_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09561_ (.A1(_02519_),
    .A2(_03699_),
    .B(_03700_),
    .C(_02798_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09562_ (.A1(_00874_),
    .A2(_01021_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09563_ (.A1(_00783_),
    .A2(_03702_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09564_ (.A1(_00796_),
    .A2(_03703_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09565_ (.A1(_03701_),
    .A2(_03704_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09566_ (.I(_02821_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09567_ (.I(_00665_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09568_ (.A1(_03707_),
    .A2(_00742_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09569_ (.I(_00510_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09570_ (.I(_00790_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09571_ (.I(_03710_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09572_ (.A1(_03706_),
    .A2(_03708_),
    .B(_03709_),
    .C(_03711_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09573_ (.A1(_00781_),
    .A2(_00731_),
    .A3(_00590_),
    .A4(_00907_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09574_ (.I(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09575_ (.A1(_00874_),
    .A2(_00890_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09576_ (.A1(_00731_),
    .A2(_03715_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09577_ (.A1(_00495_),
    .A2(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09578_ (.A1(_03705_),
    .A2(_03712_),
    .A3(_03714_),
    .A4(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09579_ (.I(_00784_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09580_ (.I(_03719_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09581_ (.A1(_00786_),
    .A2(_03707_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09582_ (.A1(_03720_),
    .A2(_00732_),
    .B(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09583_ (.A1(net26),
    .A2(_03718_),
    .B(_02999_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09584_ (.A1(_03718_),
    .A2(_03722_),
    .B(_03723_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09585_ (.I(_02529_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09586_ (.A1(_00506_),
    .A2(_00525_),
    .A3(_03724_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09587_ (.A1(net24),
    .A2(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09588_ (.A1(_05723_),
    .A2(_03725_),
    .B(_03726_),
    .C(_02926_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09589_ (.A1(_00501_),
    .A2(_02512_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(_00885_),
    .A2(_01790_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09591_ (.A1(_02562_),
    .A2(_03728_),
    .B(_00941_),
    .C(_00886_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09592_ (.A1(_00773_),
    .A2(_00906_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09593_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09594_ (.A1(_00698_),
    .A2(_03731_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09595_ (.A1(_00510_),
    .A2(_02557_),
    .A3(_00863_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(_03732_),
    .A2(_03733_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09597_ (.A1(_00649_),
    .A2(_02516_),
    .A3(_03734_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09598_ (.A1(_02560_),
    .A2(_03729_),
    .B(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09599_ (.I0(net25),
    .I1(_03727_),
    .S(_03736_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09600_ (.A1(_00857_),
    .A2(_03737_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09601_ (.I(_03738_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09602_ (.I(_00975_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09603_ (.A1(_02514_),
    .A2(_00731_),
    .A3(_00592_),
    .A4(_00907_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09604_ (.A1(_00981_),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09605_ (.I(_02525_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09606_ (.A1(_00764_),
    .A2(_00597_),
    .A3(_03716_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09607_ (.A1(_03742_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09608_ (.A1(\as2650.cycle[9] ),
    .A2(_03739_),
    .A3(_03741_),
    .B(_03744_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09609_ (.A1(_00609_),
    .A2(_02544_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09610_ (.I(_03746_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09611_ (.A1(_00647_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .B(_00497_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09612_ (.A1(_00764_),
    .A2(_01782_),
    .A3(_02552_),
    .B(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09613_ (.A1(_00597_),
    .A2(_01786_),
    .A3(_03731_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09614_ (.A1(_02515_),
    .A2(_00703_),
    .B(_03749_),
    .C(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09615_ (.A1(_00615_),
    .A2(_02544_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09616_ (.A1(_00815_),
    .A2(_03752_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09617_ (.A1(_05733_),
    .A2(_00485_),
    .A3(_00605_),
    .A4(_02511_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09618_ (.A1(_03753_),
    .A2(_03754_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09619_ (.A1(_00661_),
    .A2(_03747_),
    .B(_03751_),
    .C(_03755_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09620_ (.I(_00602_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09621_ (.I(_02533_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09622_ (.A1(_00789_),
    .A2(_02529_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09623_ (.A1(_03757_),
    .A2(_00946_),
    .A3(_03758_),
    .A4(_03759_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09624_ (.A1(_02550_),
    .A2(_02568_),
    .A3(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09625_ (.A1(_00875_),
    .A2(_00595_),
    .A3(_01189_),
    .A4(_02797_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09626_ (.A1(_01809_),
    .A2(_02538_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09627_ (.A1(_00613_),
    .A2(_03731_),
    .B(_03762_),
    .C(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09628_ (.A1(_03745_),
    .A2(_03756_),
    .A3(_03761_),
    .A4(_03764_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09629_ (.A1(_00455_),
    .A2(_00485_),
    .A3(_00676_),
    .A4(_02512_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09630_ (.A1(_02358_),
    .A2(_02531_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09631_ (.A1(_02515_),
    .A2(_01782_),
    .A3(_02557_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09632_ (.A1(_00689_),
    .A2(_00672_),
    .A3(_01790_),
    .A4(_02797_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09633_ (.A1(_00816_),
    .A2(_00960_),
    .A3(_03724_),
    .B(_03769_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09634_ (.A1(_00636_),
    .A2(_03768_),
    .B(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09635_ (.I(_02553_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09636_ (.A1(_00691_),
    .A2(_02572_),
    .A3(_02511_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09637_ (.A1(_00781_),
    .A2(_02529_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09638_ (.A1(_00478_),
    .A2(_02790_),
    .A3(_00960_),
    .A4(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09639_ (.A1(_05727_),
    .A2(_00944_),
    .A3(_00688_),
    .A4(_02554_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09640_ (.A1(_02527_),
    .A2(_03776_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09641_ (.A1(_03772_),
    .A2(_03773_),
    .A3(_03775_),
    .A4(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09642_ (.A1(_03767_),
    .A2(_03771_),
    .A3(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09643_ (.A1(_03766_),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09644_ (.A1(_03765_),
    .A2(_03780_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09645_ (.I(_03781_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09646_ (.I(_03782_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09647_ (.I(net93),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09648_ (.I(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09649_ (.I(_03785_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09650_ (.I(_00569_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09651_ (.A1(_03787_),
    .A2(_02587_),
    .B(_02596_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09652_ (.I(_03788_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09653_ (.I(_00560_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09654_ (.I(_03790_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09655_ (.I(_00978_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09656_ (.A1(_01091_),
    .A2(_01086_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09657_ (.A1(_01115_),
    .A2(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09658_ (.A1(_03792_),
    .A2(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09659_ (.I(_01436_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09660_ (.A1(_03796_),
    .A2(_03793_),
    .B(_02864_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09661_ (.I(_00557_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09662_ (.A1(\as2650.cycle[10] ),
    .A2(\as2650.cycle[2] ),
    .B(_00758_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09663_ (.I(_03799_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09664_ (.A1(_03798_),
    .A2(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09665_ (.A1(_00750_),
    .A2(_00574_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09666_ (.A1(_00748_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09667_ (.I(net99),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09668_ (.A1(_03795_),
    .A2(_03797_),
    .A3(_03801_),
    .B1(_03803_),
    .B2(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(_03791_),
    .A2(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09670_ (.I(_01026_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09671_ (.A1(_03807_),
    .A2(_01098_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09672_ (.A1(_02863_),
    .A2(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09673_ (.A1(_01819_),
    .A2(_01117_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09674_ (.A1(_00570_),
    .A2(_02821_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09675_ (.A1(_00562_),
    .A2(_03809_),
    .B1(_03810_),
    .B2(_00547_),
    .C(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_03806_),
    .A2(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09677_ (.I(_00634_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09678_ (.A1(_00642_),
    .A2(_00596_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09679_ (.I(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09680_ (.A1(_03814_),
    .A2(_02812_),
    .A3(_03816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09681_ (.I(_03817_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09682_ (.I(_00868_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09683_ (.A1(_03804_),
    .A2(_00869_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09684_ (.A1(_03819_),
    .A2(_03810_),
    .B(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09685_ (.A1(_00671_),
    .A2(_00616_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09686_ (.I(net99),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09687_ (.I(_00706_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09688_ (.A1(_03823_),
    .A2(_03824_),
    .B1(_00722_),
    .B2(_01117_),
    .C(_00993_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09689_ (.A1(_03823_),
    .A2(_01785_),
    .B(_03825_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09690_ (.A1(_03786_),
    .A2(_03822_),
    .B(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09691_ (.A1(_01820_),
    .A2(_02852_),
    .B1(_00719_),
    .B2(_03827_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09692_ (.A1(_03818_),
    .A2(_03821_),
    .B(_03828_),
    .C(_00791_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09693_ (.A1(_02671_),
    .A2(_03711_),
    .B(_00785_),
    .C(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09694_ (.A1(_03813_),
    .A2(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09695_ (.A1(_03786_),
    .A2(_03789_),
    .B1(_03831_),
    .B2(_02598_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09696_ (.I(_03781_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09697_ (.I(_03833_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09698_ (.A1(_03804_),
    .A2(_03834_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09699_ (.I(_00754_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09700_ (.A1(_03783_),
    .A2(_03832_),
    .B(_03835_),
    .C(_03836_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09701_ (.I(_03782_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09702_ (.I(net92),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09703_ (.I(_03788_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09704_ (.I(_00759_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09705_ (.I(_02864_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09706_ (.A1(net92),
    .A2(_01208_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09707_ (.A1(_03786_),
    .A2(_03841_),
    .A3(_03842_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09708_ (.I(_00546_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09709_ (.A1(_03784_),
    .A2(_01115_),
    .B(_03842_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09710_ (.A1(_03844_),
    .A2(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09711_ (.I(_02784_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09712_ (.I(_01211_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09713_ (.A1(_01210_),
    .A2(_01229_),
    .A3(_03794_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09714_ (.A1(_00978_),
    .A2(_03849_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09715_ (.A1(_03848_),
    .A2(_03792_),
    .B(_03850_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09716_ (.A1(_00563_),
    .A2(_01025_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09717_ (.I(_03852_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09718_ (.A1(_01115_),
    .A2(_01097_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09719_ (.A1(_02981_),
    .A2(_01199_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09720_ (.A1(_03854_),
    .A2(_03855_),
    .B(_03807_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09721_ (.A1(_03854_),
    .A2(_03855_),
    .B(_03856_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09722_ (.A1(_03848_),
    .A2(_03853_),
    .B(_03857_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09723_ (.A1(_03800_),
    .A2(_03851_),
    .B1(_03858_),
    .B2(_00579_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09724_ (.I(net31),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09725_ (.A1(_03860_),
    .A2(_03804_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09726_ (.I(_03790_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09727_ (.A1(_00748_),
    .A2(_03859_),
    .B1(_03861_),
    .B2(_03803_),
    .C(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09728_ (.A1(_03843_),
    .A2(_03846_),
    .B(_03847_),
    .C(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09729_ (.I(_02519_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09730_ (.A1(_03784_),
    .A2(_01116_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09731_ (.A1(_03866_),
    .A2(_03842_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09732_ (.I0(_03860_),
    .I1(_03867_),
    .S(_02961_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09733_ (.I(_00667_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09734_ (.A1(_00634_),
    .A2(_00779_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09735_ (.I(_03870_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09736_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09737_ (.A1(_03869_),
    .A2(_03872_),
    .B(_01835_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09738_ (.I(_02814_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09739_ (.I(_00616_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09740_ (.A1(_00673_),
    .A2(_03875_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09741_ (.I(_00722_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09742_ (.A1(_02865_),
    .A2(_03877_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09743_ (.A1(_00564_),
    .A2(_00610_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09744_ (.I(_03879_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09745_ (.A1(_03860_),
    .A2(_03880_),
    .B1(_03861_),
    .B2(_00741_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09746_ (.A1(_03874_),
    .A2(_03876_),
    .A3(_03878_),
    .A4(_03881_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09747_ (.A1(_03818_),
    .A2(_03868_),
    .B(_03873_),
    .C(_03882_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09748_ (.I(_00840_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09749_ (.A1(_01836_),
    .A2(_03865_),
    .B1(_03883_),
    .B2(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09750_ (.A1(_03864_),
    .A2(_03885_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09751_ (.A1(_03840_),
    .A2(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09752_ (.A1(_03838_),
    .A2(_03839_),
    .B(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09753_ (.A1(_03860_),
    .A2(_03834_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09754_ (.A1(_03837_),
    .A2(_03888_),
    .B(_03889_),
    .C(_03836_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09755_ (.I(net32),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09756_ (.I(net57),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09757_ (.I(_03891_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09758_ (.I(_00783_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09759_ (.I(_03893_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09760_ (.I(_03822_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09761_ (.A1(_00824_),
    .A2(_02569_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09762_ (.I(_03896_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09763_ (.A1(_03895_),
    .A2(_03897_),
    .B(_03892_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09764_ (.I(_00673_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09765_ (.I(_00993_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09766_ (.I(_03900_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09767_ (.I(_03901_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09768_ (.A1(_00563_),
    .A2(_00654_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09769_ (.I(_03903_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09770_ (.A1(net31),
    .A2(net99),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09771_ (.A1(_03890_),
    .A2(_03905_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09772_ (.I(_00655_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09773_ (.I(_03907_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09774_ (.I(_01785_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _09775_ (.A1(_02867_),
    .A2(_03904_),
    .B1(_03906_),
    .B2(_03908_),
    .C1(_03909_),
    .C2(_03890_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09776_ (.I(_02961_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09777_ (.I(_00833_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09778_ (.A1(_01855_),
    .A2(_01251_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09779_ (.A1(net56),
    .A2(_01208_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09780_ (.A1(net93),
    .A2(net8),
    .A3(_03842_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09781_ (.A1(_03914_),
    .A2(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09782_ (.A1(_03913_),
    .A2(_03916_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09783_ (.I(_03817_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09784_ (.A1(_03912_),
    .A2(_03917_),
    .B(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09785_ (.A1(_03890_),
    .A2(_03911_),
    .B(_03919_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09786_ (.A1(_03899_),
    .A2(_03902_),
    .A3(_03910_),
    .B(_03920_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09787_ (.I(_03884_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09788_ (.I(_01436_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09789_ (.I(net10),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09790_ (.I(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09791_ (.A1(_01209_),
    .A2(_01228_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09792_ (.A1(_01209_),
    .A2(_01228_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09793_ (.A1(_03794_),
    .A2(_03926_),
    .B(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09794_ (.A1(_03925_),
    .A2(_01274_),
    .A3(_03928_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09795_ (.A1(_02866_),
    .A2(_03923_),
    .B(_03800_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09796_ (.A1(_03923_),
    .A2(_03929_),
    .B(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09797_ (.I(_01026_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09798_ (.A1(_01209_),
    .A2(_01200_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09799_ (.A1(_03854_),
    .A2(_03855_),
    .B(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09800_ (.A1(_03925_),
    .A2(_01269_),
    .A3(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09801_ (.I(_02866_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09802_ (.A1(_03936_),
    .A2(_03807_),
    .B(_00578_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09803_ (.A1(_03932_),
    .A2(_03935_),
    .B(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09804_ (.A1(_03931_),
    .A2(_03938_),
    .B(_03798_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09805_ (.A1(_00574_),
    .A2(_00578_),
    .B(_00557_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09806_ (.A1(_03940_),
    .A2(_03906_),
    .B(_00547_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09807_ (.A1(_03891_),
    .A2(net10),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09808_ (.A1(_03914_),
    .A2(_03845_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09809_ (.A1(_03942_),
    .A2(_03943_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09810_ (.A1(_03939_),
    .A2(_03941_),
    .B1(_03944_),
    .B2(_03844_),
    .C(_03811_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09811_ (.A1(_03894_),
    .A2(_03898_),
    .B1(_03921_),
    .B2(_03922_),
    .C(_03945_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09812_ (.A1(_03892_),
    .A2(_03789_),
    .B1(_03946_),
    .B2(_02597_),
    .C(_03782_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09813_ (.A1(_03890_),
    .A2(_03837_),
    .B(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09814_ (.A1(_02926_),
    .A2(_03948_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09815_ (.I(_03834_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09816_ (.I(_00748_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09817_ (.A1(_03936_),
    .A2(_01275_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09818_ (.A1(_01252_),
    .A2(_01274_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(_03928_),
    .A2(_03952_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09820_ (.A1(_02871_),
    .A2(_01367_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09821_ (.A1(_03951_),
    .A2(_03953_),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09822_ (.A1(_03951_),
    .A2(_03954_),
    .A3(_03953_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09823_ (.I(_03923_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09824_ (.A1(_03955_),
    .A2(_03956_),
    .B(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09825_ (.I(_03739_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09826_ (.A1(_02873_),
    .A2(_03792_),
    .B(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09827_ (.I(_03853_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09828_ (.A1(_01348_),
    .A2(_01362_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09829_ (.A1(_01263_),
    .A2(net81),
    .B(_03925_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09830_ (.A1(_03924_),
    .A2(_01263_),
    .A3(net81),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09831_ (.A1(_03934_),
    .A2(_03963_),
    .B(_03964_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09832_ (.A1(_03962_),
    .A2(_03965_),
    .B(_03932_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09833_ (.A1(_03962_),
    .A2(_03965_),
    .B(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09834_ (.A1(_02873_),
    .A2(_03961_),
    .B(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09835_ (.I(_00579_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09836_ (.A1(_03958_),
    .A2(_03960_),
    .B1(_03968_),
    .B2(_03969_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09837_ (.I(net98),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09838_ (.A1(net32),
    .A2(net31),
    .A3(net99),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09839_ (.A1(_03971_),
    .A2(_03972_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09840_ (.I(_03803_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09841_ (.I(_03790_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09842_ (.A1(_03950_),
    .A2(_03970_),
    .B1(_03973_),
    .B2(_03974_),
    .C(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09843_ (.I(net58),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(_03977_),
    .A2(_01348_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09845_ (.A1(_01866_),
    .A2(_02870_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09846_ (.A1(_03978_),
    .A2(_03979_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_01854_),
    .A2(_01251_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_03913_),
    .A2(_03943_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(_03981_),
    .A2(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09850_ (.A1(_03980_),
    .A2(_03983_),
    .B(_03791_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09851_ (.A1(_03980_),
    .A2(_03983_),
    .B(_03984_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09852_ (.A1(_03840_),
    .A2(_03847_),
    .A3(_03976_),
    .A4(_03985_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09853_ (.I(_03710_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09854_ (.A1(_03987_),
    .A2(_03706_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09855_ (.A1(_00742_),
    .A2(_03973_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09856_ (.I(_03879_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09857_ (.A1(_02873_),
    .A2(_00723_),
    .B1(_03990_),
    .B2(net98),
    .C(_03816_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09858_ (.I(_00868_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09859_ (.I(_03992_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(_03814_),
    .A2(_03816_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09861_ (.I(_03994_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09862_ (.I(_00867_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09863_ (.I(_03996_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09864_ (.A1(_03942_),
    .A2(_03916_),
    .B(_03981_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09865_ (.A1(_03980_),
    .A2(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09866_ (.A1(_03997_),
    .A2(_03999_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09867_ (.A1(net98),
    .A2(_03993_),
    .B(_03995_),
    .C(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09868_ (.A1(_03989_),
    .A2(_03991_),
    .B(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09869_ (.I(_03977_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09870_ (.I(_03822_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09871_ (.A1(_04004_),
    .A2(_03896_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09872_ (.I(_04005_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(_04003_),
    .A2(_04006_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09874_ (.A1(_03988_),
    .A2(_04002_),
    .B(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09875_ (.A1(_00570_),
    .A2(_02596_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09876_ (.A1(_04008_),
    .A2(_04009_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09877_ (.A1(_01867_),
    .A2(_03839_),
    .B(_03986_),
    .C(_04010_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09878_ (.I(_03833_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(net98),
    .A2(_04012_),
    .B(_02999_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09880_ (.A1(_03949_),
    .A2(_04011_),
    .B(_04013_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09881_ (.I(_00759_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09882_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09883_ (.A1(_02869_),
    .A2(_01367_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09884_ (.A1(_01252_),
    .A2(_01274_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09885_ (.A1(_01347_),
    .A2(_01366_),
    .B1(_03928_),
    .B2(_03952_),
    .C(_04017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09886_ (.A1(_04016_),
    .A2(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09887_ (.A1(_02976_),
    .A2(_01428_),
    .A3(_04019_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09888_ (.I(_03800_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09889_ (.A1(_02876_),
    .A2(_03957_),
    .B(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09890_ (.A1(_03957_),
    .A2(_04020_),
    .B(_04022_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09891_ (.A1(_02869_),
    .A2(_01361_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09892_ (.A1(_02869_),
    .A2(_01361_),
    .B1(_03934_),
    .B2(_03963_),
    .C(_03964_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09893_ (.A1(_04024_),
    .A2(_04025_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09894_ (.A1(_01409_),
    .A2(_01403_),
    .A3(_04026_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09895_ (.I(_00578_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09896_ (.A1(_03961_),
    .A2(_04027_),
    .B(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09897_ (.A1(_02976_),
    .A2(_03961_),
    .B(_04029_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09898_ (.I(_00557_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09899_ (.A1(_04023_),
    .A2(_04030_),
    .B(_04031_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09900_ (.I(_03940_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09901_ (.I(net34),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09902_ (.A1(_03971_),
    .A2(_03972_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09903_ (.A1(_04034_),
    .A2(_04035_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_00547_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09905_ (.A1(_04033_),
    .A2(_04036_),
    .B(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09906_ (.A1(_01878_),
    .A2(_01406_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09907_ (.A1(_03978_),
    .A2(_03983_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09908_ (.A1(_03979_),
    .A2(_04040_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09909_ (.A1(_04039_),
    .A2(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09910_ (.I(_03811_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09911_ (.A1(_04032_),
    .A2(_04038_),
    .B1(_04042_),
    .B2(_00548_),
    .C(_04043_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09912_ (.A1(_00784_),
    .A2(_00704_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09913_ (.I(_04045_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09914_ (.I(_01878_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _09915_ (.A1(_02875_),
    .A2(_03904_),
    .B1(_04036_),
    .B2(_00881_),
    .C1(_03909_),
    .C2(_04034_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09916_ (.A1(_03977_),
    .A2(_01348_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09917_ (.A1(_03978_),
    .A2(_03998_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09918_ (.A1(_04049_),
    .A2(_04050_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09919_ (.A1(_04039_),
    .A2(_04051_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09920_ (.A1(_00553_),
    .A2(_04052_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09921_ (.A1(_04034_),
    .A2(_03911_),
    .B(_04053_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09922_ (.A1(_03816_),
    .A2(_04048_),
    .B1(_04054_),
    .B2(_03995_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09923_ (.I(_03896_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09924_ (.A1(_04047_),
    .A2(_04006_),
    .B1(_04055_),
    .B2(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09925_ (.A1(_01880_),
    .A2(_03789_),
    .B1(_04046_),
    .B2(_04057_),
    .C(_03833_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09926_ (.A1(_04015_),
    .A2(_04044_),
    .B(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09927_ (.I(_00829_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09928_ (.A1(_04034_),
    .A2(_03837_),
    .B(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09929_ (.A1(_04059_),
    .A2(_04061_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09930_ (.I(net35),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09931_ (.I(_01192_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09932_ (.A1(_01407_),
    .A2(_01403_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09933_ (.A1(_01407_),
    .A2(_01403_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09934_ (.A1(_04024_),
    .A2(_04064_),
    .A3(_04025_),
    .B(_04065_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09935_ (.A1(_01501_),
    .A2(_01509_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09936_ (.A1(_04066_),
    .A2(_04067_),
    .B(_03853_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09937_ (.A1(_04066_),
    .A2(_04067_),
    .B(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09938_ (.A1(_02584_),
    .A2(_03932_),
    .B(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09939_ (.A1(_01406_),
    .A2(_01427_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09940_ (.A1(_01407_),
    .A2(_01427_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09941_ (.A1(_04016_),
    .A2(_04071_),
    .A3(_04018_),
    .B(_04072_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09942_ (.A1(_01500_),
    .A2(_01493_),
    .A3(_04073_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09943_ (.A1(_03796_),
    .A2(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09944_ (.A1(_02583_),
    .A2(_03796_),
    .B(_04075_),
    .C(_04021_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09945_ (.A1(_04063_),
    .A2(_04070_),
    .B(_04076_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09946_ (.A1(net34),
    .A2(_04035_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09947_ (.A1(net35),
    .A2(_04078_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09948_ (.A1(_03974_),
    .A2(_04079_),
    .B(_03791_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09949_ (.A1(_04031_),
    .A2(_04077_),
    .B(_04080_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09950_ (.A1(_01893_),
    .A2(_01498_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09951_ (.I(_04082_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09952_ (.A1(net60),
    .A2(net12),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09953_ (.A1(_04039_),
    .A2(_04041_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09954_ (.A1(_04084_),
    .A2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09955_ (.A1(_04083_),
    .A2(_04086_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09956_ (.A1(_03975_),
    .A2(_04087_),
    .B(_03847_),
    .C(_00760_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09957_ (.A1(_04081_),
    .A2(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09958_ (.I(_01892_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09959_ (.I(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09960_ (.A1(_02591_),
    .A2(_00723_),
    .B1(_04079_),
    .B2(_00708_),
    .C1(_03990_),
    .C2(_04062_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09961_ (.A1(_03876_),
    .A2(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09962_ (.A1(_04049_),
    .A2(_04050_),
    .B(_04039_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09963_ (.A1(_04084_),
    .A2(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09964_ (.A1(_04083_),
    .A2(_04095_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09965_ (.A1(_04062_),
    .A2(_00869_),
    .B(_03994_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09966_ (.A1(_03993_),
    .A2(_04096_),
    .B(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04093_),
    .A2(_04098_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09968_ (.A1(_01894_),
    .A2(_04005_),
    .B1(_04099_),
    .B2(_03897_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09969_ (.A1(_04091_),
    .A2(_03788_),
    .B1(_04046_),
    .B2(_04100_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09970_ (.A1(_04089_),
    .A2(_04101_),
    .B(_03782_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09971_ (.A1(_04062_),
    .A2(_04012_),
    .B(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09972_ (.A1(_02926_),
    .A2(_04103_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09973_ (.I(_03862_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09974_ (.I(_01571_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09975_ (.I(_04105_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09976_ (.I(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09977_ (.A1(_04106_),
    .A2(_01596_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09978_ (.A1(_01498_),
    .A2(_01492_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09979_ (.A1(_01499_),
    .A2(_01492_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09980_ (.A1(_04073_),
    .A2(_04109_),
    .B(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09981_ (.A1(_04108_),
    .A2(_04111_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09982_ (.A1(_03923_),
    .A2(_04112_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09983_ (.A1(_04107_),
    .A2(_03796_),
    .B(_04113_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09984_ (.A1(_04106_),
    .A2(_01591_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09985_ (.A1(_04107_),
    .A2(_01592_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09986_ (.A1(_04115_),
    .A2(_04116_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09987_ (.A1(_01499_),
    .A2(_01508_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09988_ (.A1(_01499_),
    .A2(_01508_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09989_ (.A1(_04066_),
    .A2(_04118_),
    .B(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09990_ (.A1(_04117_),
    .A2(_04120_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09991_ (.A1(_03807_),
    .A2(_04121_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09992_ (.A1(_04107_),
    .A2(_03932_),
    .B(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09993_ (.I(_01192_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09994_ (.A1(_03739_),
    .A2(_04114_),
    .B1(_04123_),
    .B2(_04124_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09995_ (.I(net36),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09996_ (.A1(_04062_),
    .A2(_04078_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09997_ (.A1(_04126_),
    .A2(_04127_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09998_ (.A1(_03798_),
    .A2(_04125_),
    .B1(_04128_),
    .B2(_03940_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09999_ (.A1(_04085_),
    .A2(_04083_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10000_ (.A1(net61),
    .A2(net1),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10001_ (.A1(_04091_),
    .A2(_01501_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10002_ (.A1(_04084_),
    .A2(_04131_),
    .B(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10003_ (.A1(net62),
    .A2(_01571_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10004_ (.I(_04134_),
    .Z(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10005_ (.A1(_04130_),
    .A2(_04133_),
    .B(_04135_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10006_ (.A1(_04135_),
    .A2(_04130_),
    .A3(_04133_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10007_ (.A1(_03791_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10008_ (.I(_03811_),
    .Z(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10009_ (.A1(_04104_),
    .A2(_04129_),
    .B1(_04136_),
    .B2(_04138_),
    .C(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10010_ (.A1(_04084_),
    .A2(_04131_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10011_ (.A1(_01892_),
    .A2(net1),
    .B(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10012_ (.A1(_04094_),
    .A2(_04082_),
    .B(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10013_ (.A1(_04135_),
    .A2(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10014_ (.A1(_03997_),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10015_ (.I(_00552_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10016_ (.A1(_04126_),
    .A2(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10017_ (.I(_00610_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10018_ (.I(_04148_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10019_ (.A1(_04149_),
    .A2(_04128_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10020_ (.A1(_02877_),
    .A2(_03904_),
    .B1(_03909_),
    .B2(_04126_),
    .C(_03876_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10021_ (.A1(_03995_),
    .A2(_04145_),
    .A3(_04147_),
    .B1(_04150_),
    .B2(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10022_ (.I(_00570_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10023_ (.A1(_01906_),
    .A2(_04006_),
    .B1(_04152_),
    .B2(_04056_),
    .C(_04153_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04140_),
    .A2(_04154_),
    .B(_03840_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10025_ (.A1(_01906_),
    .A2(_03789_),
    .B(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10026_ (.A1(_04126_),
    .A2(_03834_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10027_ (.A1(_03837_),
    .A2(_04156_),
    .B(_04157_),
    .C(_03836_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_03788_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10029_ (.A1(_01573_),
    .A2(_01597_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10030_ (.A1(_04108_),
    .A2(_04111_),
    .B(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10031_ (.A1(_02960_),
    .A2(_01692_),
    .A3(_04160_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10032_ (.A1(_03957_),
    .A2(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10033_ (.A1(_00835_),
    .A2(_03792_),
    .B(_03959_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10034_ (.A1(_04117_),
    .A2(_04120_),
    .B(_04115_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10035_ (.A1(_02960_),
    .A2(_01687_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10036_ (.A1(_04164_),
    .A2(_04165_),
    .B(_03853_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10037_ (.A1(_04164_),
    .A2(_04165_),
    .B(_04166_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10038_ (.I(_01192_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10039_ (.A1(_00835_),
    .A2(_03961_),
    .B(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10040_ (.A1(_04162_),
    .A2(_04163_),
    .B1(_04167_),
    .B2(_04169_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10041_ (.I(net37),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10042_ (.A1(net36),
    .A2(net35),
    .A3(_04078_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10043_ (.A1(_04171_),
    .A2(_04172_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10044_ (.A1(_04033_),
    .A2(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10045_ (.A1(_03950_),
    .A2(_04170_),
    .B(_04174_),
    .C(_04104_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10046_ (.A1(net63),
    .A2(net2),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10047_ (.A1(_01905_),
    .A2(_01571_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10048_ (.A1(_04177_),
    .A2(_04136_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10049_ (.A1(_04176_),
    .A2(_04178_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10050_ (.A1(_04037_),
    .A2(_04179_),
    .B(_04043_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10051_ (.I(_03897_),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10052_ (.I(_00551_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10053_ (.A1(_04182_),
    .A2(_00722_),
    .B1(_03880_),
    .B2(_04171_),
    .C(_03900_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10054_ (.A1(_03908_),
    .A2(_04173_),
    .B(_04183_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10055_ (.A1(_01919_),
    .A2(_03895_),
    .B(_04184_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10056_ (.A1(_04135_),
    .A2(_04143_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10057_ (.A1(_04177_),
    .A2(_04186_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10058_ (.A1(_04176_),
    .A2(_04187_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10059_ (.A1(_00869_),
    .A2(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10060_ (.A1(_04171_),
    .A2(_03997_),
    .B(_03918_),
    .C(_04189_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10061_ (.A1(_00838_),
    .A2(_04185_),
    .B(_04190_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10062_ (.A1(_01919_),
    .A2(_04181_),
    .B1(_04191_),
    .B2(_00826_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10063_ (.I(_00785_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10064_ (.A1(_04175_),
    .A2(_04180_),
    .B1(_04192_),
    .B2(_04193_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10065_ (.I(_02596_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10066_ (.A1(_01919_),
    .A2(_04158_),
    .B1(_04194_),
    .B2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10067_ (.A1(_04171_),
    .A2(_04012_),
    .B(_02999_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10068_ (.A1(_03949_),
    .A2(_04196_),
    .B(_04197_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10069_ (.I(\as2650.addr_buff[0] ),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10070_ (.A1(_00549_),
    .A2(_01691_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10071_ (.A1(_04108_),
    .A2(_04111_),
    .B(_04199_),
    .C(_04159_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10072_ (.A1(_00831_),
    .A2(_01691_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10073_ (.A1(_00978_),
    .A2(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10074_ (.A1(_04200_),
    .A2(_04202_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10075_ (.A1(_04198_),
    .A2(_04203_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10076_ (.I(_04198_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10077_ (.A1(_00831_),
    .A2(_01686_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10078_ (.A1(_04117_),
    .A2(_04120_),
    .B(_04206_),
    .C(_04115_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10079_ (.A1(_00550_),
    .A2(_01686_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10080_ (.A1(_03852_),
    .A2(_04208_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10081_ (.A1(_04207_),
    .A2(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10082_ (.A1(_04205_),
    .A2(_04210_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10083_ (.A1(_04021_),
    .A2(_04204_),
    .B1(_04211_),
    .B2(_04028_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10084_ (.I(net38),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10085_ (.I(net37),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10086_ (.A1(_04214_),
    .A2(_04172_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10087_ (.A1(_04213_),
    .A2(_04215_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10088_ (.A1(_03950_),
    .A2(_04212_),
    .B1(_04216_),
    .B2(_03974_),
    .C(_03975_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10089_ (.A1(net91),
    .A2(_01572_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10090_ (.A1(_04134_),
    .A2(_04176_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10091_ (.A1(_04142_),
    .A2(_04219_),
    .B(_04177_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10092_ (.A1(_01918_),
    .A2(_01572_),
    .B(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10093_ (.A1(_04085_),
    .A2(_04083_),
    .A3(_04219_),
    .B(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10094_ (.A1(_04218_),
    .A2(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10095_ (.A1(_04218_),
    .A2(_04222_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10096_ (.A1(_03975_),
    .A2(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10097_ (.A1(_04223_),
    .A2(_04225_),
    .B(_04139_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10098_ (.A1(_00881_),
    .A2(_04216_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10099_ (.A1(_04205_),
    .A2(_03904_),
    .B1(_03909_),
    .B2(_04213_),
    .C(_03876_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10100_ (.A1(_04094_),
    .A2(_04082_),
    .A3(_04219_),
    .B(_04221_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10101_ (.A1(_04218_),
    .A2(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10102_ (.A1(_00553_),
    .A2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10103_ (.A1(_04213_),
    .A2(_03911_),
    .B(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10104_ (.A1(_04227_),
    .A2(_04228_),
    .B1(_04232_),
    .B2(_03995_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10105_ (.A1(_02214_),
    .A2(_04006_),
    .B1(_04233_),
    .B2(_04056_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10106_ (.A1(_04217_),
    .A2(_04226_),
    .B1(_04234_),
    .B2(_04193_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10107_ (.I(_02597_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10108_ (.A1(_02214_),
    .A2(_04158_),
    .B1(_04235_),
    .B2(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10109_ (.I(_02998_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10110_ (.A1(_04213_),
    .A2(_04012_),
    .B(_04238_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10111_ (.A1(_03949_),
    .A2(_04237_),
    .B(_04239_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10112_ (.I(net39),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10113_ (.A1(net38),
    .A2(_04215_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10114_ (.A1(_04240_),
    .A2(_04241_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10115_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10116_ (.A1(_04210_),
    .A2(_04243_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10117_ (.I(_04198_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10118_ (.I(\as2650.addr_buff[1] ),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10119_ (.A1(_04245_),
    .A2(_04210_),
    .B(_04246_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10120_ (.A1(_04244_),
    .A2(_04247_),
    .B(_04168_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10121_ (.A1(_04203_),
    .A2(_04243_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10122_ (.A1(_04245_),
    .A2(_04203_),
    .B(_04246_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10123_ (.A1(_04249_),
    .A2(_04250_),
    .B(_03959_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10124_ (.A1(_04248_),
    .A2(_04251_),
    .B(_04031_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10125_ (.A1(_03974_),
    .A2(_04242_),
    .B(_04252_),
    .C(_04104_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10126_ (.I(net65),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10127_ (.I(_04254_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10128_ (.I(_04105_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10129_ (.A1(_04255_),
    .A2(_04256_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10130_ (.I(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(_02212_),
    .A2(_01575_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10132_ (.A1(_04259_),
    .A2(_04223_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10133_ (.A1(_04258_),
    .A2(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10134_ (.A1(_04037_),
    .A2(_04261_),
    .B(_04139_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10135_ (.A1(_00708_),
    .A2(_04242_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10136_ (.I(\as2650.addr_buff[1] ),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10137_ (.A1(_04264_),
    .A2(_03877_),
    .B1(_03880_),
    .B2(_04240_),
    .C(_03900_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10138_ (.A1(_04255_),
    .A2(_03872_),
    .B1(_04263_),
    .B2(_04265_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(_04218_),
    .A2(_04229_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10140_ (.A1(_04259_),
    .A2(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10141_ (.A1(_04258_),
    .A2(_04268_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10142_ (.I(_00868_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(_04240_),
    .A2(_04270_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10144_ (.A1(_03819_),
    .A2(_04269_),
    .B(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10145_ (.A1(_00674_),
    .A2(_04266_),
    .B1(_04272_),
    .B2(_03918_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10146_ (.A1(_03987_),
    .A2(_04273_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10147_ (.A1(_02226_),
    .A2(_04181_),
    .B(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10148_ (.A1(_04253_),
    .A2(_04262_),
    .B1(_04275_),
    .B2(_04193_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10149_ (.A1(_02226_),
    .A2(_04158_),
    .B1(_04276_),
    .B2(_04236_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10150_ (.I(_03833_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10151_ (.A1(_04240_),
    .A2(_04278_),
    .B(_04238_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10152_ (.A1(_03949_),
    .A2(_04277_),
    .B(_04279_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10153_ (.A1(net66),
    .A2(_04105_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10154_ (.I(_04280_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10155_ (.A1(_02225_),
    .A2(net91),
    .B(_04256_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10156_ (.A1(_04267_),
    .A2(_04257_),
    .B(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10157_ (.A1(_04281_),
    .A2(_04283_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10158_ (.A1(_03997_),
    .A2(_04284_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10159_ (.A1(net97),
    .A2(_04146_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10160_ (.I(_03871_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10161_ (.I(\as2650.addr_buff[2] ),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10162_ (.A1(net39),
    .A2(net38),
    .A3(_04215_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10163_ (.A1(net97),
    .A2(_04289_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10164_ (.I(_00707_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10165_ (.I(net97),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10166_ (.A1(_04288_),
    .A2(_03877_),
    .B1(_04290_),
    .B2(_04291_),
    .C1(_03990_),
    .C2(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10167_ (.I(_01190_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10168_ (.A1(_02234_),
    .A2(_04287_),
    .B1(_04293_),
    .B2(_04294_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10169_ (.I(_00673_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10170_ (.I(_04296_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10171_ (.A1(_03818_),
    .A2(_04285_),
    .A3(_04286_),
    .B1(_04295_),
    .B2(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10172_ (.A1(_02234_),
    .A2(_03988_),
    .B1(_04298_),
    .B2(_00792_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10173_ (.A1(_04288_),
    .A2(_04243_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10174_ (.A1(_04207_),
    .A2(_04209_),
    .A3(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(_04288_),
    .A2(_04244_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10176_ (.A1(_04301_),
    .A2(_04302_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10177_ (.A1(_04200_),
    .A2(_04202_),
    .A3(_04300_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10178_ (.A1(_04288_),
    .A2(_04249_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10179_ (.A1(_04304_),
    .A2(_04305_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10180_ (.A1(_03969_),
    .A2(_04303_),
    .B1(_04306_),
    .B2(_04021_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(_04033_),
    .A2(_04290_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10182_ (.A1(_03950_),
    .A2(_04307_),
    .B(_04308_),
    .C(_04104_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10183_ (.A1(_04223_),
    .A2(_04258_),
    .B(_04282_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10184_ (.A1(_04281_),
    .A2(_04310_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10185_ (.A1(_04037_),
    .A2(_04311_),
    .B(_04043_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10186_ (.A1(_04193_),
    .A2(_04299_),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10187_ (.A1(_02234_),
    .A2(_03839_),
    .B1(_04313_),
    .B2(_04236_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10188_ (.A1(net97),
    .A2(_04278_),
    .B(_04238_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10189_ (.A1(_03783_),
    .A2(_04314_),
    .B(_04315_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10190_ (.A1(net67),
    .A2(_01572_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10191_ (.A1(_02232_),
    .A2(_04256_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10192_ (.A1(_04281_),
    .A2(_04310_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10193_ (.A1(_04317_),
    .A2(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10194_ (.A1(_04316_),
    .A2(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10195_ (.I(\as2650.addr_buff[3] ),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10196_ (.I(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10197_ (.A1(_04322_),
    .A2(_04301_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10198_ (.A1(_04322_),
    .A2(_04304_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10199_ (.A1(_04168_),
    .A2(_04323_),
    .B1(_04324_),
    .B2(_03959_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10200_ (.I(net41),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10201_ (.A1(_04292_),
    .A2(_04289_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10202_ (.A1(_04326_),
    .A2(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10203_ (.A1(_04031_),
    .A2(_04325_),
    .B1(_04328_),
    .B2(_04033_),
    .C(_03844_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10204_ (.A1(_00548_),
    .A2(_04320_),
    .B(_04329_),
    .C(_04043_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10205_ (.I(_00718_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10206_ (.I(_04331_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10207_ (.I(\as2650.addr_buff[3] ),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10208_ (.A1(_04333_),
    .A2(_03877_),
    .B1(_03880_),
    .B2(_04326_),
    .C(_02804_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10209_ (.A1(_03908_),
    .A2(_04328_),
    .B(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10210_ (.A1(_02240_),
    .A2(_03895_),
    .B(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10211_ (.A1(_04281_),
    .A2(_04283_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10212_ (.A1(_04317_),
    .A2(_04337_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10213_ (.A1(_04316_),
    .A2(_04338_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10214_ (.A1(_00835_),
    .A2(_04339_),
    .B(_03918_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10215_ (.A1(_04326_),
    .A2(_03993_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10216_ (.A1(_04332_),
    .A2(_04336_),
    .B1(_04340_),
    .B2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10217_ (.A1(_02240_),
    .A2(_04153_),
    .A3(_04181_),
    .B1(_04342_),
    .B2(_00464_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10218_ (.I(_00760_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10219_ (.A1(_04330_),
    .A2(_04343_),
    .B(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10220_ (.A1(_02240_),
    .A2(_04158_),
    .B(_04345_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10221_ (.A1(_04326_),
    .A2(_04278_),
    .B(_04238_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10222_ (.A1(_03783_),
    .A2(_04346_),
    .B(_04347_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10223_ (.I(_03893_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10224_ (.A1(_02246_),
    .A2(_04056_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10225_ (.I(_02245_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10226_ (.A1(net41),
    .A2(_04327_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10227_ (.A1(net96),
    .A2(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10228_ (.A1(_00742_),
    .A2(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10229_ (.I(\as2650.addr_buff[4] ),
    .Z(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10230_ (.I(_03900_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10231_ (.A1(_04354_),
    .A2(_00723_),
    .B1(_03990_),
    .B2(net96),
    .C(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10232_ (.A1(_04350_),
    .A2(_04287_),
    .B1(_04353_),
    .B2(_04356_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10233_ (.A1(net68),
    .A2(_01573_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10234_ (.A1(_04280_),
    .A2(_04316_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10235_ (.A1(_04317_),
    .A2(_04282_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10236_ (.A1(_02238_),
    .A2(_01573_),
    .B(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10237_ (.A1(_04267_),
    .A2(_04257_),
    .A3(_04359_),
    .B(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10238_ (.A1(_04358_),
    .A2(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10239_ (.A1(net96),
    .A2(_03993_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10240_ (.A1(_00870_),
    .A2(_04363_),
    .B(_04364_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10241_ (.A1(_00675_),
    .A2(_04357_),
    .B1(_04365_),
    .B2(_03818_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10242_ (.I(_03884_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10243_ (.A1(_04223_),
    .A2(_04258_),
    .A3(_04359_),
    .B(_04361_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10244_ (.A1(_04358_),
    .A2(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10245_ (.I(\as2650.addr_buff[4] ),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10246_ (.A1(_04322_),
    .A2(_04301_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10247_ (.A1(_04370_),
    .A2(_04371_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10248_ (.A1(_04321_),
    .A2(_04304_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10249_ (.A1(_04370_),
    .A2(_04373_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10250_ (.A1(_04124_),
    .A2(_04372_),
    .B1(_04374_),
    .B2(_03739_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10251_ (.A1(_03803_),
    .A2(_04352_),
    .B(_03862_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10252_ (.A1(_03798_),
    .A2(_04375_),
    .B(_04376_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10253_ (.A1(_03844_),
    .A2(_04369_),
    .B(_04377_),
    .C(_04139_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10254_ (.A1(_04348_),
    .A2(_04349_),
    .B1(_04366_),
    .B2(_04367_),
    .C(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10255_ (.A1(_02246_),
    .A2(_03839_),
    .B1(_04379_),
    .B2(_04236_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _10256_ (.I(_00828_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10257_ (.A1(net96),
    .A2(_04278_),
    .B(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10258_ (.A1(_03783_),
    .A2(_04380_),
    .B(_04382_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10259_ (.A1(_02568_),
    .A2(_03773_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10260_ (.A1(_02538_),
    .A2(_04383_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10261_ (.A1(_03767_),
    .A2(_03777_),
    .A3(_04384_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10262_ (.A1(_00739_),
    .A2(_02794_),
    .A3(_03732_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10263_ (.I(_00867_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10264_ (.A1(_04387_),
    .A2(_03790_),
    .B(_00749_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10265_ (.A1(_00858_),
    .A2(_04388_),
    .B(_03740_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10266_ (.A1(_03771_),
    .A2(_04386_),
    .A3(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10267_ (.A1(_03745_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10268_ (.A1(_02556_),
    .A2(_03775_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10269_ (.A1(_00694_),
    .A2(_03768_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10270_ (.A1(_00883_),
    .A2(_02370_),
    .A3(_03703_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10271_ (.I(_00518_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10272_ (.I(_00841_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10273_ (.A1(_04395_),
    .A2(_04396_),
    .A3(_01784_),
    .A4(_02370_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10274_ (.A1(_04393_),
    .A2(_03661_),
    .A3(_04394_),
    .A4(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10275_ (.A1(_00750_),
    .A2(_00575_),
    .A3(_03741_),
    .B(_03755_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10276_ (.A1(_03735_),
    .A2(_04392_),
    .A3(_04398_),
    .A4(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10277_ (.A1(_04385_),
    .A2(_04391_),
    .A3(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10278_ (.A1(_03766_),
    .A2(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10279_ (.I(_00791_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10280_ (.I(_00526_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10281_ (.I(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10282_ (.I(_00668_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10283_ (.A1(net85),
    .A2(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10284_ (.A1(_03706_),
    .A2(_03709_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10285_ (.A1(_04405_),
    .A2(_04407_),
    .B(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10286_ (.A1(net95),
    .A2(_00623_),
    .B(_00589_),
    .C(_03847_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10287_ (.A1(net95),
    .A2(_00849_),
    .A3(_04181_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10288_ (.A1(_04403_),
    .A2(_04409_),
    .B(_04410_),
    .C(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10289_ (.A1(_04015_),
    .A2(_04412_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10290_ (.A1(net95),
    .A2(_04402_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10291_ (.A1(_04402_),
    .A2(_04413_),
    .B(_04414_),
    .C(_03836_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10292_ (.I(net94),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10293_ (.A1(_00765_),
    .A2(_00462_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10294_ (.A1(_03757_),
    .A2(_02812_),
    .A3(_02960_),
    .A4(_00780_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _10295_ (.A1(_02569_),
    .A2(_00486_),
    .A3(_03822_),
    .B1(_04417_),
    .B2(_00787_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10296_ (.A1(_00839_),
    .A2(_00516_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10297_ (.I(_04419_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10298_ (.A1(_04420_),
    .A2(_00606_),
    .A3(_00612_),
    .A4(_03747_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10299_ (.A1(_00642_),
    .A2(_00604_),
    .A3(_01021_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10300_ (.A1(_00714_),
    .A2(_00659_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _10301_ (.A1(_04420_),
    .A2(_00716_),
    .A3(_00660_),
    .B1(_04422_),
    .B2(_04423_),
    .B3(_00657_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10302_ (.A1(_04149_),
    .A2(_02545_),
    .A3(_04424_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10303_ (.A1(_00953_),
    .A2(_00698_),
    .A3(_00520_),
    .A4(_03752_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10304_ (.A1(_03754_),
    .A2(_03749_),
    .A3(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10305_ (.I(_02568_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10306_ (.A1(_01783_),
    .A2(_04393_),
    .A3(_03734_),
    .A4(_03744_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10307_ (.A1(_02555_),
    .A2(_04428_),
    .A3(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10308_ (.A1(_04425_),
    .A2(_04427_),
    .A3(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10309_ (.A1(_04416_),
    .A2(_04418_),
    .B(_04421_),
    .C(_04431_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10310_ (.A1(_03780_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10311_ (.A1(_00766_),
    .A2(_00758_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10312_ (.A1(net94),
    .A2(_04153_),
    .A3(_00778_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10313_ (.I(_00655_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10314_ (.I(_00628_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10315_ (.A1(_00715_),
    .A2(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10316_ (.A1(_00847_),
    .A2(_00970_),
    .A3(_04436_),
    .B1(_03903_),
    .B2(_04438_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10317_ (.A1(net94),
    .A2(_04439_),
    .B(_04296_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10318_ (.A1(_03911_),
    .A2(_04331_),
    .B(_03710_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10319_ (.A1(net94),
    .A2(_00824_),
    .A3(_03709_),
    .A4(_00729_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10320_ (.A1(_04440_),
    .A2(_04441_),
    .B(_04442_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10321_ (.A1(_03719_),
    .A2(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10322_ (.A1(_00970_),
    .A2(_04435_),
    .B(_04444_),
    .C(_02545_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10323_ (.A1(_04434_),
    .A2(_04445_),
    .B(_04433_),
    .C(_02598_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10324_ (.I(_00754_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10325_ (.A1(_04415_),
    .A2(_04433_),
    .B(_04446_),
    .C(_04447_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10326_ (.A1(_00714_),
    .A2(_00862_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10327_ (.A1(_00843_),
    .A2(_04448_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10328_ (.A1(_00732_),
    .A2(_00598_),
    .B(_03715_),
    .C(_00779_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10329_ (.A1(_00569_),
    .A2(_01020_),
    .A3(_03136_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10330_ (.A1(_00981_),
    .A2(_03799_),
    .A3(_03714_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10331_ (.A1(_00677_),
    .A2(_04450_),
    .B(_04451_),
    .C(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10332_ (.A1(_00527_),
    .A2(_00639_),
    .A3(_02545_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10333_ (.A1(_00546_),
    .A2(_03714_),
    .B(_04454_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10334_ (.A1(_03704_),
    .A2(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10335_ (.A1(_00883_),
    .A2(_00718_),
    .A3(_02785_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10336_ (.A1(_04453_),
    .A2(_04456_),
    .A3(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10337_ (.I(_01190_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10338_ (.I(_03824_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10339_ (.A1(_00519_),
    .A2(_00706_),
    .A3(_00611_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10340_ (.A1(_04460_),
    .A2(_04423_),
    .A3(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10341_ (.A1(_00840_),
    .A2(_00719_),
    .A3(_04459_),
    .A4(_04462_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10342_ (.A1(_02959_),
    .A2(_04449_),
    .B(_04458_),
    .C(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10343_ (.I(_04464_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10344_ (.I0(_03841_),
    .I1(_04205_),
    .S(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10345_ (.I(_04466_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10346_ (.I(_04465_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10347_ (.I(_04464_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10348_ (.A1(_04264_),
    .A2(_04468_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10349_ (.A1(_02981_),
    .A2(_04467_),
    .B(_04469_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10350_ (.I(\as2650.addr_buff[2] ),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10351_ (.I(_04464_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_04470_),
    .A2(_04471_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10353_ (.A1(_03925_),
    .A2(_04467_),
    .B(_04472_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(_04333_),
    .A2(_04471_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10355_ (.A1(_01349_),
    .A2(_04467_),
    .B(_04473_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_04354_),
    .A2(_04471_),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10357_ (.A1(_02976_),
    .A2(_04467_),
    .B(_04474_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10358_ (.A1(_01024_),
    .A2(_04471_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10359_ (.A1(_02584_),
    .A2(_04468_),
    .B(_04475_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10360_ (.I(_01023_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10361_ (.A1(_04476_),
    .A2(_04465_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10362_ (.A1(_04107_),
    .A2(_04468_),
    .B(_04477_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10363_ (.A1(_00565_),
    .A2(_04465_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10364_ (.A1(_00870_),
    .A2(_04468_),
    .B(_04478_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10365_ (.A1(\as2650.last_intr ),
    .A2(_04195_),
    .B(_04381_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10366_ (.A1(_00647_),
    .A2(_04195_),
    .B(_04479_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10367_ (.I(_00902_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10368_ (.I(_04480_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10369_ (.A1(_04481_),
    .A2(_04060_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10370_ (.A1(_01016_),
    .A2(_04482_),
    .B(_02560_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10371_ (.A1(_00765_),
    .A2(_00816_),
    .A3(_03702_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10372_ (.A1(_00546_),
    .A2(_03740_),
    .B(_03743_),
    .C(_04483_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10373_ (.A1(_00746_),
    .A2(_04063_),
    .B(_03862_),
    .C(_03740_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10374_ (.A1(_00817_),
    .A2(_03724_),
    .B(_01783_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10375_ (.A1(_02856_),
    .A2(_02560_),
    .B(_03753_),
    .C(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10376_ (.A1(_03751_),
    .A2(_04484_),
    .A3(_04485_),
    .A4(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10377_ (.A1(_01024_),
    .A2(_04015_),
    .B(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10378_ (.A1(_01082_),
    .A2(_04488_),
    .B(_04489_),
    .C(_04447_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10379_ (.A1(_04476_),
    .A2(_04015_),
    .B(_04488_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10380_ (.A1(_01084_),
    .A2(_04488_),
    .B(_04490_),
    .C(_04447_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10381_ (.I(_00998_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10382_ (.A1(_00962_),
    .A2(_01056_),
    .B(_00806_),
    .C(_01055_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10383_ (.A1(_03869_),
    .A2(_02790_),
    .A3(_04492_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10384_ (.A1(_04491_),
    .A2(_04493_),
    .B(_00883_),
    .C(_01017_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10385_ (.I(_04494_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10386_ (.I(_04495_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10387_ (.I(_02812_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_04497_),
    .A2(_02864_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10389_ (.A1(_01137_),
    .A2(_02570_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(_04498_),
    .A2(_04499_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10391_ (.A1(_04496_),
    .A2(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10392_ (.A1(_01043_),
    .A2(_04496_),
    .B(_04501_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10393_ (.I(_04494_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10394_ (.I(_02364_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10395_ (.A1(_01239_),
    .A2(_02959_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10396_ (.A1(_04503_),
    .A2(_02981_),
    .B(_04504_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10397_ (.A1(_04502_),
    .A2(_04505_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10398_ (.A1(_01163_),
    .A2(_04496_),
    .B(_04506_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10399_ (.I(_02569_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10400_ (.I(_04507_),
    .Z(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10401_ (.I(_00538_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10402_ (.A1(_04509_),
    .A2(_02867_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10403_ (.A1(_01847_),
    .A2(_04508_),
    .B(_04510_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10404_ (.I0(_04511_),
    .I1(\as2650.holding_reg[2] ),
    .S(_04502_),
    .Z(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10405_ (.I(_04512_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10406_ (.A1(_02133_),
    .A2(_04406_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10407_ (.A1(_02581_),
    .A2(_01349_),
    .B(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10408_ (.I0(_04514_),
    .I1(\as2650.holding_reg[3] ),
    .S(_04502_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10409_ (.I(_04515_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10410_ (.A1(_02156_),
    .A2(_02588_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10411_ (.I(_02876_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10412_ (.A1(_02823_),
    .A2(_04517_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10413_ (.A1(_04516_),
    .A2(_04518_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10414_ (.I0(_04519_),
    .I1(\as2650.holding_reg[4] ),
    .S(_04495_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10415_ (.I(_04520_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10416_ (.A1(_01496_),
    .A2(_04507_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10417_ (.A1(_00539_),
    .A2(_02583_),
    .B(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10418_ (.A1(_04502_),
    .A2(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10419_ (.A1(_01515_),
    .A2(_04496_),
    .B(_04523_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10420_ (.I(_02877_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10421_ (.A1(_02823_),
    .A2(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10422_ (.A1(_03672_),
    .A2(_02581_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10423_ (.A1(_04525_),
    .A2(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10424_ (.I0(_04527_),
    .I1(\as2650.holding_reg[6] ),
    .S(_04495_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10425_ (.I(_04528_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10426_ (.A1(_02822_),
    .A2(_04146_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10427_ (.A1(_04529_),
    .A2(_02365_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10428_ (.I0(_04530_),
    .I1(\as2650.holding_reg[7] ),
    .S(_04495_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10429_ (.I(_04531_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10430_ (.A1(_00902_),
    .A2(_00720_),
    .A3(_00729_),
    .A4(_04529_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10431_ (.A1(_00766_),
    .A2(_04532_),
    .B(_00733_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10432_ (.I(_04533_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10433_ (.I(_00775_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10434_ (.A1(_00767_),
    .A2(_03841_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10435_ (.A1(_05711_),
    .A2(_04534_),
    .B1(_04535_),
    .B2(_04536_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10436_ (.I(_02865_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10437_ (.A1(_00767_),
    .A2(_04537_),
    .B(_04416_),
    .C(_04533_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10438_ (.A1(_01932_),
    .A2(_04534_),
    .B(_04538_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10439_ (.A1(_00788_),
    .A2(_04534_),
    .B1(_00776_),
    .B2(_02868_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10440_ (.I(_04539_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10441_ (.A1(_00767_),
    .A2(_02591_),
    .B1(_00721_),
    .B2(_04416_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10442_ (.A1(_00679_),
    .A2(_04535_),
    .B1(_04540_),
    .B2(_04534_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10443_ (.A1(_00805_),
    .A2(_04533_),
    .B1(_00776_),
    .B2(_04524_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10444_ (.I(_04541_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10445_ (.A1(_00804_),
    .A2(_04533_),
    .B1(_00776_),
    .B2(_00836_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10446_ (.I(_04542_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10447_ (.A1(_00816_),
    .A2(_00960_),
    .A3(_03724_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10448_ (.A1(_00885_),
    .A2(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10449_ (.A1(_03748_),
    .A2(_04544_),
    .B(_00755_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10450_ (.A1(_02515_),
    .A2(_00598_),
    .A3(_04422_),
    .A4(_04461_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10451_ (.A1(_02561_),
    .A2(_04545_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(_03741_),
    .A2(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10453_ (.A1(_02517_),
    .A2(_03750_),
    .A3(_04543_),
    .A4(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10454_ (.A1(_03757_),
    .A2(_00946_),
    .A3(_03758_),
    .A4(_03759_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10455_ (.A1(_03772_),
    .A2(_04549_),
    .A3(_03775_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10456_ (.A1(_04420_),
    .A2(_00716_),
    .A3(_00660_),
    .A4(_03747_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10457_ (.A1(_00657_),
    .A2(_03747_),
    .A3(_04422_),
    .A4(_04423_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10458_ (.A1(_04419_),
    .A2(_00606_),
    .A3(_00612_),
    .A4(_03746_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10459_ (.A1(_00796_),
    .A2(_02558_),
    .B(_03753_),
    .C(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10460_ (.A1(_04419_),
    .A2(_03903_),
    .A3(_03815_),
    .A4(_03730_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10461_ (.I(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10462_ (.A1(_02550_),
    .A2(_04552_),
    .A3(_04554_),
    .A4(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10463_ (.A1(_02525_),
    .A2(_03748_),
    .A3(_03769_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10464_ (.A1(_04550_),
    .A2(_04551_),
    .A3(_04557_),
    .A4(_04558_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10465_ (.A1(_04385_),
    .A2(_04484_),
    .A3(_04548_),
    .A4(_04559_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10466_ (.I(_04560_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10467_ (.I(_04561_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10468_ (.I(_04562_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10469_ (.I(_04009_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10470_ (.I(_02578_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10471_ (.A1(_00825_),
    .A2(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10472_ (.I(_02783_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10473_ (.A1(\as2650.stack[7][0] ),
    .A2(_01964_),
    .B1(_02048_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10474_ (.I(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10475_ (.A1(\as2650.stack[4][0] ),
    .A2(_02004_),
    .B1(_02001_),
    .B2(\as2650.stack[5][0] ),
    .C(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10476_ (.I(_01801_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10477_ (.A1(\as2650.stack[0][0] ),
    .A2(_04571_),
    .B1(_01984_),
    .B2(\as2650.stack[2][0] ),
    .C1(_02001_),
    .C2(\as2650.stack[1][0] ),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10478_ (.A1(\as2650.stack[3][0] ),
    .A2(_02041_),
    .B(_01955_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10479_ (.A1(_01996_),
    .A2(_04570_),
    .B1(_04572_),
    .B2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10480_ (.A1(\as2650.stack[8][0] ),
    .A2(_02044_),
    .B1(_02051_),
    .B2(\as2650.stack[9][0] ),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10481_ (.A1(\as2650.stack[11][0] ),
    .A2(_02041_),
    .B1(_02071_),
    .B2(\as2650.stack[10][0] ),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10482_ (.A1(_02934_),
    .A2(_04575_),
    .A3(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10483_ (.A1(\as2650.stack[15][0] ),
    .A2(_02040_),
    .B1(_02048_),
    .B2(\as2650.stack[14][0] ),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10484_ (.I(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10485_ (.A1(\as2650.stack[12][0] ),
    .A2(_02004_),
    .B1(_02051_),
    .B2(\as2650.stack[13][0] ),
    .C(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10486_ (.A1(_01996_),
    .A2(_04580_),
    .B(_01951_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10487_ (.A1(_02008_),
    .A2(_04574_),
    .B1(_04577_),
    .B2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10488_ (.A1(_03784_),
    .A2(_00671_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10489_ (.A1(_00454_),
    .A2(_04583_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10490_ (.A1(_02670_),
    .A2(_00454_),
    .B(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10491_ (.I0(_03785_),
    .I1(_04583_),
    .S(_05733_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10492_ (.I0(_04585_),
    .I1(_04586_),
    .S(_05736_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10493_ (.A1(_03785_),
    .A2(_00552_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10494_ (.A1(_04182_),
    .A2(_03810_),
    .B(_04588_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10495_ (.A1(_04396_),
    .A2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10496_ (.I(_03870_),
    .Z(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(_01117_),
    .A2(_00656_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10498_ (.A1(_04245_),
    .A2(_03907_),
    .B(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10499_ (.A1(_02670_),
    .A2(_04591_),
    .B1(_04593_),
    .B2(_04437_),
    .C(_02586_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10500_ (.I(_00715_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10501_ (.A1(_00539_),
    .A2(_04587_),
    .B1(_04590_),
    .B2(_04594_),
    .C(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10502_ (.A1(_05805_),
    .A2(_00656_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10503_ (.A1(_02863_),
    .A2(_04597_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10504_ (.I(_01190_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10505_ (.A1(_01820_),
    .A2(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10506_ (.A1(_04294_),
    .A2(_04598_),
    .B(_04600_),
    .C(_00739_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_01820_),
    .A2(_03869_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10508_ (.A1(_00674_),
    .A2(_04602_),
    .B(_00825_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10509_ (.A1(_03896_),
    .A2(_04589_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10510_ (.A1(_04297_),
    .A2(_04596_),
    .A3(_04601_),
    .B1(_04603_),
    .B2(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10511_ (.A1(_03786_),
    .A2(_04566_),
    .B1(_04567_),
    .B2(_04582_),
    .C(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10512_ (.I(_01809_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10513_ (.A1(_04607_),
    .A2(_04009_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10514_ (.I(_04560_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10515_ (.A1(_04564_),
    .A2(_04606_),
    .B1(_04608_),
    .B2(_02671_),
    .C(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10516_ (.A1(_02671_),
    .A2(_04563_),
    .B(_04610_),
    .C(_04447_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10517_ (.I(_04608_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10518_ (.A1(_03838_),
    .A2(_03785_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10519_ (.A1(_03996_),
    .A2(_03867_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10520_ (.A1(_01835_),
    .A2(_04270_),
    .B(_04613_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10521_ (.I(_00842_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10522_ (.A1(_03848_),
    .A2(_04460_),
    .B(_00728_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10523_ (.A1(_04246_),
    .A2(_04291_),
    .B(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10524_ (.A1(_03872_),
    .A2(_04612_),
    .B1(_04614_),
    .B2(_04615_),
    .C(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10525_ (.I(_00457_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10526_ (.A1(_01818_),
    .A2(_00489_),
    .B(_01834_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(_01819_),
    .A2(_03814_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10528_ (.A1(_03838_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10529_ (.A1(_04620_),
    .A2(_04622_),
    .B(_00458_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10530_ (.A1(_04619_),
    .A2(_04612_),
    .B(_04623_),
    .C(_00668_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10531_ (.I(_00520_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10532_ (.A1(_04508_),
    .A2(_04618_),
    .B(_04624_),
    .C(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10533_ (.I(_04599_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10534_ (.I(_04612_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10535_ (.I(_04459_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10536_ (.I(_00707_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10537_ (.A1(net8),
    .A2(_05805_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10538_ (.A1(_02980_),
    .A2(_05796_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10539_ (.A1(_04631_),
    .A2(_04632_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10540_ (.A1(_04631_),
    .A2(_04632_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_04633_),
    .A2(_04634_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10542_ (.I(_03824_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10543_ (.A1(_03848_),
    .A2(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10544_ (.A1(_04630_),
    .A2(_04635_),
    .B(_04637_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10545_ (.A1(_04629_),
    .A2(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10546_ (.A1(_04627_),
    .A2(_04628_),
    .B(_04639_),
    .C(_00848_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10547_ (.A1(_04332_),
    .A2(_04626_),
    .A3(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10548_ (.A1(_04508_),
    .A2(_04628_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10549_ (.I(_04296_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10550_ (.A1(_00540_),
    .A2(_04614_),
    .B(_04642_),
    .C(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10551_ (.A1(_04403_),
    .A2(_04641_),
    .A3(_04644_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10552_ (.A1(_00790_),
    .A2(_00878_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10553_ (.I(_04646_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10554_ (.A1(\as2650.stack[7][1] ),
    .A2(_01963_),
    .B1(_02047_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10555_ (.I(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10556_ (.A1(\as2650.stack[4][1] ),
    .A2(_02043_),
    .B1(_02000_),
    .B2(\as2650.stack[5][1] ),
    .C(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10557_ (.A1(\as2650.stack[0][1] ),
    .A2(_02043_),
    .B1(_02048_),
    .B2(\as2650.stack[2][1] ),
    .C1(_02000_),
    .C2(\as2650.stack[1][1] ),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10558_ (.A1(\as2650.stack[3][1] ),
    .A2(_02040_),
    .B(_01954_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10559_ (.A1(_01987_),
    .A2(_04650_),
    .B1(_04651_),
    .B2(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10560_ (.A1(\as2650.stack[8][1] ),
    .A2(_01977_),
    .B1(_01980_),
    .B2(\as2650.stack[9][1] ),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10561_ (.A1(\as2650.stack[11][1] ),
    .A2(_02040_),
    .B1(_02070_),
    .B2(\as2650.stack[10][1] ),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10562_ (.A1(_02951_),
    .A2(_04654_),
    .A3(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10563_ (.A1(\as2650.stack[15][1] ),
    .A2(_01945_),
    .B1(_02047_),
    .B2(\as2650.stack[14][1] ),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10564_ (.I(_04657_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10565_ (.A1(\as2650.stack[12][1] ),
    .A2(_02043_),
    .B1(_01980_),
    .B2(\as2650.stack[13][1] ),
    .C(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10566_ (.A1(_01987_),
    .A2(_04659_),
    .B(_01950_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10567_ (.A1(_02020_),
    .A2(_04653_),
    .B1(_04656_),
    .B2(_04660_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10568_ (.A1(_03710_),
    .A2(_02578_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10569_ (.I(_04662_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10570_ (.A1(_04647_),
    .A2(_04628_),
    .B1(_04661_),
    .B2(_04663_),
    .C(_04046_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10571_ (.A1(_04611_),
    .A2(_04612_),
    .B1(_04645_),
    .B2(_04664_),
    .C(_04609_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10572_ (.I(_00795_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10573_ (.I(_04666_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10574_ (.A1(_01836_),
    .A2(_04563_),
    .B(_04665_),
    .C(_04667_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10575_ (.I(_04560_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10576_ (.I(_04668_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10577_ (.I(_04669_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10578_ (.I(_00842_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10579_ (.A1(_01855_),
    .A2(_02961_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10580_ (.A1(_03912_),
    .A2(_03917_),
    .B(_04672_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10581_ (.A1(_01854_),
    .A2(_03838_),
    .A3(net55),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10582_ (.I(_04674_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10583_ (.A1(_01835_),
    .A2(_02670_),
    .B(_03892_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10584_ (.A1(_04675_),
    .A2(_04676_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10585_ (.A1(_04470_),
    .A2(_00880_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10586_ (.A1(_03936_),
    .A2(_04636_),
    .B(_04437_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10587_ (.A1(_04004_),
    .A2(_04677_),
    .B1(_04678_),
    .B2(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10588_ (.A1(_04671_),
    .A2(_04673_),
    .B(_04680_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10589_ (.I(_02958_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10590_ (.I(_00457_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10591_ (.A1(_01854_),
    .A2(_04620_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10592_ (.A1(_01855_),
    .A2(_04620_),
    .B(_00457_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10593_ (.A1(_04683_),
    .A2(_04677_),
    .B1(_04684_),
    .B2(_04685_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10594_ (.A1(_04682_),
    .A2(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10595_ (.A1(_02571_),
    .A2(_04681_),
    .B(_04687_),
    .C(_04625_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10596_ (.I(_04677_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10597_ (.A1(net10),
    .A2(_05789_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10598_ (.A1(_01251_),
    .A2(_05789_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10599_ (.A1(_04690_),
    .A2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10600_ (.A1(_01208_),
    .A2(_05796_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10601_ (.A1(_04693_),
    .A2(_04634_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10602_ (.A1(_04692_),
    .A2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10603_ (.A1(_03936_),
    .A2(_04636_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10604_ (.A1(_04630_),
    .A2(_04695_),
    .B(_04696_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10605_ (.A1(_04629_),
    .A2(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10606_ (.I(_00847_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10607_ (.A1(_04627_),
    .A2(_04689_),
    .B(_04698_),
    .C(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10608_ (.A1(_04332_),
    .A2(_04688_),
    .A3(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10609_ (.A1(_02571_),
    .A2(_04689_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10610_ (.A1(_00540_),
    .A2(_04673_),
    .B(_04702_),
    .C(_04643_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10611_ (.A1(_04403_),
    .A2(_04701_),
    .A3(_04703_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10612_ (.A1(\as2650.stack[8][2] ),
    .A2(_02946_),
    .B1(_02935_),
    .B2(\as2650.stack[9][2] ),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10613_ (.A1(\as2650.stack[11][2] ),
    .A2(_02945_),
    .B1(_01969_),
    .B2(\as2650.stack[10][2] ),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10614_ (.A1(_02951_),
    .A2(_04705_),
    .A3(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10615_ (.A1(\as2650.stack[15][2] ),
    .A2(_02945_),
    .B1(_02935_),
    .B2(\as2650.stack[13][2] ),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10616_ (.A1(\as2650.stack[12][2] ),
    .A2(_02946_),
    .B1(_02948_),
    .B2(\as2650.stack[14][2] ),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10617_ (.A1(_02940_),
    .A2(_04708_),
    .A3(_04709_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10618_ (.A1(_04707_),
    .A2(_04710_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10619_ (.A1(\as2650.stack[7][2] ),
    .A2(_01974_),
    .B1(_02948_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10620_ (.A1(\as2650.stack[4][2] ),
    .A2(_01977_),
    .B1(_01980_),
    .B2(\as2650.stack[5][2] ),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10621_ (.A1(_01955_),
    .A2(_04712_),
    .A3(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10622_ (.A1(\as2650.stack[0][2] ),
    .A2(_01977_),
    .B1(_01960_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10623_ (.A1(\as2650.stack[3][2] ),
    .A2(_01974_),
    .B1(_02070_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10624_ (.A1(_02951_),
    .A2(_04715_),
    .A3(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10625_ (.A1(_02020_),
    .A2(_04714_),
    .A3(_04717_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10626_ (.A1(_01951_),
    .A2(_04711_),
    .B(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _10627_ (.I(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10628_ (.A1(_04647_),
    .A2(_04689_),
    .B1(_04720_),
    .B2(_04663_),
    .C(_04046_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10629_ (.I(_04607_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10630_ (.A1(_04722_),
    .A2(_04009_),
    .A3(_04689_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10631_ (.A1(_04704_),
    .A2(_04721_),
    .B(_04723_),
    .C(_04562_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10632_ (.A1(_03892_),
    .A2(_04670_),
    .B(_04724_),
    .C(_04667_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10633_ (.A1(_04003_),
    .A2(_04675_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10634_ (.A1(_01866_),
    .A2(_04675_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10635_ (.A1(\as2650.stack[8][3] ),
    .A2(_01978_),
    .B1(_01961_),
    .B2(\as2650.stack[9][3] ),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10636_ (.A1(\as2650.stack[11][3] ),
    .A2(_01975_),
    .B1(_02150_),
    .B2(\as2650.stack[10][3] ),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10637_ (.A1(_02032_),
    .A2(_04727_),
    .A3(_04728_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10638_ (.A1(\as2650.stack[14][3] ),
    .A2(_02150_),
    .B1(_01981_),
    .B2(\as2650.stack[13][3] ),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10639_ (.A1(\as2650.stack[15][3] ),
    .A2(_01992_),
    .B1(_01978_),
    .B2(\as2650.stack[12][3] ),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10640_ (.A1(_01956_),
    .A2(_04730_),
    .A3(_04731_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10641_ (.A1(_04729_),
    .A2(_04732_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10642_ (.A1(\as2650.stack[7][3] ),
    .A2(_01992_),
    .B1(_02150_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10643_ (.A1(\as2650.stack[4][3] ),
    .A2(_02044_),
    .B1(_01981_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10644_ (.A1(_01988_),
    .A2(_04734_),
    .A3(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10645_ (.A1(\as2650.stack[2][3] ),
    .A2(_02071_),
    .B1(_01981_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10646_ (.A1(\as2650.stack[3][3] ),
    .A2(_01992_),
    .B1(_01978_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10647_ (.A1(_02032_),
    .A2(_04737_),
    .A3(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10648_ (.A1(_02021_),
    .A2(_04736_),
    .A3(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10649_ (.A1(_01952_),
    .A2(_04733_),
    .B(_04740_),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10650_ (.I(_04741_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_01867_),
    .A2(_04182_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10652_ (.A1(_00834_),
    .A2(_03999_),
    .B(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_04615_),
    .A2(_04744_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10654_ (.A1(_04322_),
    .A2(_00741_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10655_ (.A1(_01349_),
    .A2(_00880_),
    .B(_03875_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10656_ (.A1(_04591_),
    .A2(_04725_),
    .B1(_04746_),
    .B2(_04747_),
    .C(_02364_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10657_ (.A1(_01866_),
    .A2(_04684_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(_02893_),
    .A2(_04726_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(_02958_),
    .A2(_00458_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10660_ (.A1(_04683_),
    .A2(_04749_),
    .B1(_04750_),
    .B2(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10661_ (.A1(_04745_),
    .A2(_04748_),
    .B(_04395_),
    .C(_04752_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10662_ (.A1(_00668_),
    .A2(_04744_),
    .B(_04750_),
    .C(_04296_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10663_ (.A1(net11),
    .A2(_05784_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10664_ (.A1(_04693_),
    .A2(_04634_),
    .B(_04690_),
    .C(_04691_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10665_ (.A1(_04690_),
    .A2(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10666_ (.A1(_04755_),
    .A2(_04757_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10667_ (.A1(_02872_),
    .A2(_04148_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10668_ (.A1(_04291_),
    .A2(_04758_),
    .B(_04759_),
    .C(_04459_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10669_ (.A1(_04294_),
    .A2(_04725_),
    .B(_04760_),
    .C(_04595_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10670_ (.A1(_00791_),
    .A2(_04754_),
    .A3(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10671_ (.A1(_04753_),
    .A2(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10672_ (.A1(_04647_),
    .A2(_04726_),
    .B1(_04742_),
    .B2(_04663_),
    .C(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10673_ (.A1(_04611_),
    .A2(_04725_),
    .B1(_04764_),
    .B2(_04564_),
    .C(_04609_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10674_ (.A1(_04003_),
    .A2(_04670_),
    .B(_04765_),
    .C(_04667_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10675_ (.A1(_04003_),
    .A2(_04675_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10676_ (.A1(_04047_),
    .A2(_04766_),
    .Z(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10677_ (.A1(_02875_),
    .A2(_04636_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(_01347_),
    .A2(_05784_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10679_ (.A1(_04690_),
    .A2(_04756_),
    .B(_04755_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10680_ (.A1(net12),
    .A2(_05772_),
    .Z(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10681_ (.I(_04771_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10682_ (.A1(_04769_),
    .A2(_04770_),
    .A3(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10683_ (.A1(_04769_),
    .A2(_04770_),
    .B(_04772_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10684_ (.A1(_00708_),
    .A2(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10685_ (.A1(_04773_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10686_ (.I(_02804_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10687_ (.A1(_04768_),
    .A2(_04776_),
    .B(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10688_ (.A1(_03902_),
    .A2(_04767_),
    .B(_04778_),
    .C(_00522_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _10689_ (.A1(_01878_),
    .A2(net58),
    .A3(_04684_),
    .Z(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10690_ (.A1(_01867_),
    .A2(_04684_),
    .B(_04047_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10691_ (.A1(_04780_),
    .A2(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10692_ (.I(_04767_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10693_ (.A1(_04507_),
    .A2(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10694_ (.A1(_04619_),
    .A2(_04782_),
    .B1(_04784_),
    .B2(_04751_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_04047_),
    .A2(_04182_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10696_ (.A1(_00834_),
    .A2(_04052_),
    .B(_04786_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10697_ (.A1(_04370_),
    .A2(_04460_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10698_ (.A1(_02875_),
    .A2(_03907_),
    .B(_00667_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10699_ (.A1(_04788_),
    .A2(_04789_),
    .B(_04491_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10700_ (.A1(_03872_),
    .A2(_04767_),
    .B1(_04787_),
    .B2(_04615_),
    .C(_04790_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10701_ (.A1(_04395_),
    .A2(_04785_),
    .A3(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10702_ (.A1(_04699_),
    .A2(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10703_ (.A1(_02853_),
    .A2(_04787_),
    .B(_04784_),
    .C(_04643_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10704_ (.A1(_04779_),
    .A2(_04793_),
    .B(_04794_),
    .C(_04403_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10705_ (.A1(\as2650.stack[7][4] ),
    .A2(_01965_),
    .B1(_01984_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10706_ (.I(_04796_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10707_ (.A1(\as2650.stack[4][4] ),
    .A2(_02005_),
    .B1(_02002_),
    .B2(\as2650.stack[5][4] ),
    .C(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10708_ (.A1(\as2650.stack[0][4] ),
    .A2(_01803_),
    .B1(_01970_),
    .B2(\as2650.stack[2][4] ),
    .C1(_01961_),
    .C2(\as2650.stack[1][4] ),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10709_ (.A1(\as2650.stack[3][4] ),
    .A2(_01966_),
    .B(_01988_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10710_ (.A1(_01999_),
    .A2(_04798_),
    .B1(_04799_),
    .B2(_04800_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10711_ (.A1(\as2650.stack[8][4] ),
    .A2(_02110_),
    .B1(_02067_),
    .B2(\as2650.stack[9][4] ),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10712_ (.A1(\as2650.stack[11][4] ),
    .A2(_02106_),
    .B1(_02076_),
    .B2(\as2650.stack[10][4] ),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10713_ (.A1(_02032_),
    .A2(_04802_),
    .A3(_04803_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10714_ (.A1(\as2650.stack[15][4] ),
    .A2(_02105_),
    .B1(_01984_),
    .B2(\as2650.stack[14][4] ),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10715_ (.I(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10716_ (.A1(\as2650.stack[12][4] ),
    .A2(_02005_),
    .B1(_02113_),
    .B2(\as2650.stack[13][4] ),
    .C(_04806_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10717_ (.A1(_01997_),
    .A2(_04807_),
    .B(_02021_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _10718_ (.A1(_01952_),
    .A2(_04801_),
    .B1(_04804_),
    .B2(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10719_ (.A1(_04647_),
    .A2(_04783_),
    .B1(_04809_),
    .B2(_04663_),
    .C(_04045_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10720_ (.A1(_04611_),
    .A2(_04767_),
    .B1(_04795_),
    .B2(_04810_),
    .C(_04668_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10721_ (.A1(_01880_),
    .A2(_04670_),
    .B(_04811_),
    .C(_04667_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10722_ (.I(_04562_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10723_ (.A1(_01879_),
    .A2(_03977_),
    .A3(_04674_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10724_ (.A1(_04091_),
    .A2(_04813_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10725_ (.I(_04814_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10726_ (.A1(_01406_),
    .A2(_05772_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10727_ (.A1(net1),
    .A2(_05763_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10728_ (.A1(_04816_),
    .A2(_04774_),
    .A3(_04817_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10729_ (.A1(_04816_),
    .A2(_04774_),
    .B(_04817_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10730_ (.A1(_04818_),
    .A2(_04819_),
    .B(_04460_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10731_ (.A1(_02583_),
    .A2(_04630_),
    .B(_03901_),
    .C(_04820_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10732_ (.A1(_04777_),
    .A2(_04814_),
    .B(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10733_ (.A1(_05733_),
    .A2(_00455_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10734_ (.I(_04823_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10735_ (.A1(_01894_),
    .A2(_04780_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10736_ (.A1(_04824_),
    .A2(_04814_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10737_ (.A1(_04824_),
    .A2(_04825_),
    .B(_04826_),
    .C(_04507_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10738_ (.A1(_03871_),
    .A2(_04814_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10739_ (.A1(_04091_),
    .A2(_00551_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10740_ (.A1(_00833_),
    .A2(_04096_),
    .B(_04829_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10741_ (.A1(_01092_),
    .A2(_00656_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _10742_ (.A1(_02590_),
    .A2(_00864_),
    .B1(_04830_),
    .B2(_00842_),
    .C1(_04831_),
    .C2(_00728_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10743_ (.A1(_03874_),
    .A2(_04828_),
    .A3(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10744_ (.A1(_00521_),
    .A2(_04827_),
    .A3(_04833_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10745_ (.A1(_00522_),
    .A2(_04822_),
    .B(_04834_),
    .C(_00838_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10746_ (.A1(_02580_),
    .A2(_04815_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10747_ (.A1(_03706_),
    .A2(_04830_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10748_ (.A1(_04297_),
    .A2(_04836_),
    .A3(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10749_ (.A1(_00792_),
    .A2(_04835_),
    .A3(_04838_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10750_ (.I(_04646_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10751_ (.I(_01959_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10752_ (.A1(\as2650.stack[8][5] ),
    .A2(_04571_),
    .B1(_04841_),
    .B2(\as2650.stack[9][5] ),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10753_ (.I(_01968_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10754_ (.A1(\as2650.stack[11][5] ),
    .A2(_01965_),
    .B1(_04843_),
    .B2(\as2650.stack[10][5] ),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10755_ (.A1(_02934_),
    .A2(_04842_),
    .A3(_04844_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10756_ (.A1(\as2650.stack[15][5] ),
    .A2(_01965_),
    .B1(_04843_),
    .B2(\as2650.stack[14][5] ),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10757_ (.A1(\as2650.stack[12][5] ),
    .A2(_04571_),
    .B1(_04841_),
    .B2(\as2650.stack[13][5] ),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10758_ (.A1(_02940_),
    .A2(_04846_),
    .A3(_04847_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10759_ (.A1(_04845_),
    .A2(_04848_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10760_ (.A1(\as2650.stack[4][5] ),
    .A2(_01802_),
    .B1(_04843_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10761_ (.A1(\as2650.stack[7][5] ),
    .A2(_02937_),
    .B1(_04841_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10762_ (.A1(_02940_),
    .A2(_04850_),
    .A3(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10763_ (.A1(\as2650.stack[0][5] ),
    .A2(_04571_),
    .B1(_04841_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10764_ (.A1(\as2650.stack[3][5] ),
    .A2(_02937_),
    .B1(_04843_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10765_ (.A1(_02934_),
    .A2(_04853_),
    .A3(_04854_),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10766_ (.A1(_01951_),
    .A2(_04852_),
    .A3(_04855_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10767_ (.A1(_02008_),
    .A2(_04849_),
    .B(_04856_),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10768_ (.A1(_04840_),
    .A2(_04815_),
    .B1(_04857_),
    .B2(_04662_),
    .C(_04153_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(_04839_),
    .A2(_04858_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10770_ (.A1(_03720_),
    .A2(_04815_),
    .B(_04859_),
    .C(_00761_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10771_ (.I(_04607_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10772_ (.I(_02518_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10773_ (.A1(\as2650.ivec[0] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(_04815_),
    .C(_04562_),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10774_ (.A1(_01894_),
    .A2(_04812_),
    .B1(_04860_),
    .B2(_04863_),
    .C(_00857_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_04090_),
    .A2(_04813_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10776_ (.A1(_01907_),
    .A2(_04864_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10777_ (.I(_04865_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10778_ (.A1(_04105_),
    .A2(_05834_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_01498_),
    .A2(_05763_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10780_ (.A1(_04868_),
    .A2(_04819_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10781_ (.A1(_04867_),
    .A2(_04869_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10782_ (.A1(_04149_),
    .A2(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10783_ (.A1(_02877_),
    .A2(_03908_),
    .B(_04599_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10784_ (.A1(_04355_),
    .A2(_04865_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10785_ (.A1(_04871_),
    .A2(_04872_),
    .B(_04873_),
    .C(_00787_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10786_ (.I(_04823_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(_04090_),
    .A2(_04780_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10788_ (.A1(_01906_),
    .A2(_04876_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10789_ (.A1(_04824_),
    .A2(_04877_),
    .B(_02893_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10790_ (.A1(_04875_),
    .A2(_04865_),
    .B(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(_04387_),
    .A2(_04144_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10792_ (.A1(_01907_),
    .A2(_03992_),
    .B(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10793_ (.A1(_01576_),
    .A2(_00863_),
    .B(_00892_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10794_ (.A1(_01094_),
    .A2(_03875_),
    .A3(_03907_),
    .B(_04882_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10795_ (.A1(_04591_),
    .A2(_04865_),
    .B1(_04881_),
    .B2(_04396_),
    .C(_04883_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10796_ (.A1(_00848_),
    .A2(_04879_),
    .A3(_04884_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10797_ (.A1(_04395_),
    .A2(_04874_),
    .B(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10798_ (.A1(_02959_),
    .A2(_04866_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10799_ (.A1(_03899_),
    .A2(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10800_ (.A1(_03897_),
    .A2(_04881_),
    .B1(_04888_),
    .B2(_03987_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10801_ (.I(_04646_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10802_ (.A1(_04890_),
    .A2(_04866_),
    .B(_03787_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10803_ (.A1(_04567_),
    .A2(_02921_),
    .B1(_04886_),
    .B2(_04889_),
    .C(_04891_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10804_ (.A1(_03720_),
    .A2(_04866_),
    .B(_04892_),
    .C(_00761_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10805_ (.I(_04561_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10806_ (.A1(\as2650.ivec[1] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(_04866_),
    .C(_04894_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10807_ (.A1(_01907_),
    .A2(_04812_),
    .B1(_04893_),
    .B2(_04895_),
    .C(_00857_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10808_ (.I(net63),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10809_ (.I(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10810_ (.A1(_01905_),
    .A2(_01892_),
    .A3(_04813_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10811_ (.A1(_04897_),
    .A2(_04898_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10812_ (.I(_04899_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(_03996_),
    .A2(_04188_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10814_ (.A1(_01918_),
    .A2(_04270_),
    .B(_04901_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(_02587_),
    .A2(_04900_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10816_ (.A1(_02589_),
    .A2(_04902_),
    .B(_04903_),
    .C(_04297_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10817_ (.A1(_01905_),
    .A2(_04090_),
    .A3(_04780_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10818_ (.A1(_01918_),
    .A2(_04905_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10819_ (.A1(_04824_),
    .A2(_04899_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10820_ (.A1(_04875_),
    .A2(_04906_),
    .B(_04907_),
    .C(_02570_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10821_ (.A1(_03814_),
    .A2(_00643_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_00565_),
    .A2(_03824_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10823_ (.A1(_04387_),
    .A2(_04148_),
    .B(_04910_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10824_ (.A1(_03871_),
    .A2(_04899_),
    .B1(_04911_),
    .B2(_04437_),
    .C(_00538_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10825_ (.A1(_04909_),
    .A2(_04902_),
    .B(_04912_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10826_ (.A1(_00521_),
    .A2(_04908_),
    .A3(_04913_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10827_ (.A1(_04256_),
    .A2(_05834_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10828_ (.A1(_04867_),
    .A2(_04869_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10829_ (.A1(net3),
    .A2(_05748_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10830_ (.A1(_04915_),
    .A2(_04916_),
    .B(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10831_ (.A1(_04915_),
    .A2(_04916_),
    .A3(_04917_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10832_ (.A1(_04918_),
    .A2(_04919_),
    .B(_04291_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10833_ (.A1(_03912_),
    .A2(_04436_),
    .B(_04459_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10834_ (.A1(_02804_),
    .A2(_04899_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10835_ (.A1(_04920_),
    .A2(_04921_),
    .B(_04922_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10836_ (.A1(_00848_),
    .A2(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10837_ (.A1(_00838_),
    .A2(_04914_),
    .A3(_04924_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10838_ (.A1(_00792_),
    .A2(_04904_),
    .A3(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10839_ (.A1(_04662_),
    .A2(_02956_),
    .B1(_04900_),
    .B2(_04890_),
    .C(_03787_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10840_ (.A1(_04926_),
    .A2(_04927_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10841_ (.A1(_03720_),
    .A2(_04900_),
    .B(_04928_),
    .C(_04344_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10842_ (.A1(\as2650.ivec[2] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(_04900_),
    .C(_04894_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10843_ (.I(_05700_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10844_ (.A1(_04897_),
    .A2(_04812_),
    .B1(_04929_),
    .B2(_04930_),
    .C(_04931_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10845_ (.I(net64),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10846_ (.A1(_04897_),
    .A2(_04905_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10847_ (.A1(_02213_),
    .A2(_04933_),
    .Z(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10848_ (.A1(_04896_),
    .A2(_04898_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10849_ (.A1(_02213_),
    .A2(_04935_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10850_ (.A1(_04497_),
    .A2(_04936_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10851_ (.A1(_00459_),
    .A2(_04934_),
    .B1(_04937_),
    .B2(_04751_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10852_ (.A1(_02213_),
    .A2(_03912_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10853_ (.A1(_04146_),
    .A2(_04230_),
    .B(_04939_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10854_ (.A1(_00538_),
    .A2(_02863_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10855_ (.A1(_02958_),
    .A2(_04198_),
    .A3(_00741_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10856_ (.A1(_04149_),
    .A2(_04941_),
    .B(_04942_),
    .C(_04491_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10857_ (.A1(_04287_),
    .A2(_04936_),
    .B1(_04940_),
    .B2(_04671_),
    .C(_04943_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10858_ (.A1(_04938_),
    .A2(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10859_ (.A1(_00831_),
    .A2(_05748_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10860_ (.A1(_04946_),
    .A2(_04918_),
    .B(_04148_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10861_ (.A1(_04245_),
    .A2(_04947_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10862_ (.I(_04936_),
    .Z(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10863_ (.A1(_04629_),
    .A2(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10864_ (.A1(_04627_),
    .A2(_04948_),
    .B(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10865_ (.A1(_04503_),
    .A2(_04940_),
    .B(_04937_),
    .C(_03899_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10866_ (.A1(_03884_),
    .A2(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10867_ (.A1(_00740_),
    .A2(_04945_),
    .B1(_04951_),
    .B2(_00849_),
    .C(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10868_ (.A1(_04565_),
    .A2(_04949_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10869_ (.A1(_02579_),
    .A2(_02011_),
    .B(_04955_),
    .C(_03865_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10870_ (.A1(_04348_),
    .A2(_04949_),
    .B(_04956_),
    .C(_04014_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10871_ (.I(_02518_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10872_ (.A1(\as2650.ivec[3] ),
    .A2(_04722_),
    .B1(_04958_),
    .B2(_04949_),
    .C(_04561_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10873_ (.A1(_04954_),
    .A2(_04957_),
    .B(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10874_ (.A1(_00830_),
    .A2(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10875_ (.A1(_04932_),
    .A2(_04563_),
    .B(_04961_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_02212_),
    .A2(_04935_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10877_ (.A1(_04255_),
    .A2(_04962_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10878_ (.I(_04963_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10879_ (.A1(_04254_),
    .A2(_04932_),
    .A3(_04897_),
    .A4(_04905_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10880_ (.A1(_02214_),
    .A2(_04933_),
    .B(_02226_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10881_ (.A1(_04965_),
    .A2(_04966_),
    .B(_04683_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10882_ (.A1(_00459_),
    .A2(_04964_),
    .B(_04967_),
    .C(_02580_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10883_ (.A1(_02225_),
    .A2(_00834_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10884_ (.A1(_00553_),
    .A2(_04269_),
    .B(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10885_ (.A1(_04264_),
    .A2(_04436_),
    .B(_03875_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10886_ (.A1(_04637_),
    .A2(_04971_),
    .B(_03869_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10887_ (.A1(_03895_),
    .A2(_04963_),
    .B1(_04970_),
    .B2(_04909_),
    .C(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10888_ (.A1(_00522_),
    .A2(_04968_),
    .A3(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10889_ (.A1(_04205_),
    .A2(_04947_),
    .B(_04264_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10890_ (.A1(_04946_),
    .A2(_04918_),
    .B(_00706_),
    .C(_04243_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10891_ (.A1(_04355_),
    .A2(_04975_),
    .A3(_04976_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10892_ (.A1(_03902_),
    .A2(_04963_),
    .B(_04977_),
    .C(_04625_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10893_ (.A1(_04643_),
    .A2(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10894_ (.I0(_04964_),
    .I1(_04970_),
    .S(_02822_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10895_ (.A1(_04974_),
    .A2(_04979_),
    .B1(_04980_),
    .B2(_00675_),
    .C(_00463_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10896_ (.A1(_02578_),
    .A2(_04963_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10897_ (.A1(_04565_),
    .A2(_02056_),
    .B(_04982_),
    .C(_03865_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10898_ (.A1(_04348_),
    .A2(_04964_),
    .B(_04983_),
    .C(_04014_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10899_ (.A1(\as2650.ivec[4] ),
    .A2(_04607_),
    .B1(_04958_),
    .B2(_04964_),
    .C(_04561_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_04981_),
    .A2(_04984_),
    .B(_04985_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10901_ (.A1(_04060_),
    .A2(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10902_ (.A1(_04255_),
    .A2(_04563_),
    .B(_04987_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10903_ (.I(_02232_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10904_ (.A1(\as2650.addr_buff[2] ),
    .A2(_04976_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10905_ (.A1(_04470_),
    .A2(_04976_),
    .B(_04629_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10906_ (.A1(_02225_),
    .A2(_02212_),
    .A3(_04935_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10907_ (.A1(_02233_),
    .A2(_04991_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10908_ (.I(_04992_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10909_ (.A1(_04989_),
    .A2(_04990_),
    .B1(_04993_),
    .B2(_04627_),
    .C(_04699_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10910_ (.A1(_04270_),
    .A2(_04284_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10911_ (.A1(_04988_),
    .A2(_03819_),
    .B(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_04470_),
    .A2(_00864_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10913_ (.A1(_00850_),
    .A2(_04696_),
    .B1(_04992_),
    .B2(_04004_),
    .C(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10914_ (.A1(_04671_),
    .A2(_04996_),
    .B(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10915_ (.A1(_02233_),
    .A2(_04965_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10916_ (.A1(_04875_),
    .A2(_04993_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10917_ (.A1(_04875_),
    .A2(_05000_),
    .B(_05001_),
    .C(_04509_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10918_ (.A1(_02853_),
    .A2(_04999_),
    .B(_05002_),
    .C(_04625_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10919_ (.A1(_00721_),
    .A2(_04994_),
    .A3(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10920_ (.A1(_02589_),
    .A2(_04993_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10921_ (.A1(_00540_),
    .A2(_04996_),
    .B(_05005_),
    .C(_00675_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10922_ (.A1(_04367_),
    .A2(_05004_),
    .A3(_05006_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10923_ (.A1(_04988_),
    .A2(_04991_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10924_ (.A1(_02579_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10925_ (.I(_03865_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10926_ (.A1(_02579_),
    .A2(_02096_),
    .B(_05009_),
    .C(_05010_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10927_ (.A1(_00571_),
    .A2(_04993_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10928_ (.A1(_00761_),
    .A2(_05007_),
    .A3(_05011_),
    .A4(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10929_ (.A1(\as2650.ivec[5] ),
    .A2(_04861_),
    .B1(_04862_),
    .B2(_05008_),
    .C(_04894_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10930_ (.A1(_04988_),
    .A2(_04669_),
    .B1(_05013_),
    .B2(_05014_),
    .C(_04931_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10931_ (.I(_02239_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10932_ (.A1(_04988_),
    .A2(_04991_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10933_ (.A1(_02239_),
    .A2(_05016_),
    .Z(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10934_ (.I(_05017_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10935_ (.A1(_03992_),
    .A2(_04339_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10936_ (.A1(_05015_),
    .A2(_03819_),
    .B(_05019_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(_04333_),
    .A2(_04436_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10938_ (.A1(_05021_),
    .A2(_04759_),
    .B(_00850_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10939_ (.A1(_04671_),
    .A2(_05020_),
    .B1(_05017_),
    .B2(_04287_),
    .C(_05022_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10940_ (.A1(net67),
    .A2(_02232_),
    .A3(_04965_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10941_ (.A1(_02233_),
    .A2(_04965_),
    .B(_02239_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10942_ (.A1(_05024_),
    .A2(_05025_),
    .B(_04683_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10943_ (.A1(_04619_),
    .A2(_05017_),
    .B(_05026_),
    .C(_04682_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10944_ (.A1(_02853_),
    .A2(_05023_),
    .B(_05027_),
    .C(_00740_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(_02587_),
    .A2(_05018_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10946_ (.A1(_02822_),
    .A2(_05020_),
    .B(_04331_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10947_ (.A1(\as2650.addr_buff[3] ),
    .A2(_04989_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10948_ (.A1(_03901_),
    .A2(_05031_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10949_ (.A1(_04333_),
    .A2(_04989_),
    .B(_05032_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10950_ (.A1(_04777_),
    .A2(_05017_),
    .B(_00521_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10951_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05033_),
    .B2(_05034_),
    .C(_00825_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10952_ (.A1(_05028_),
    .A2(_05035_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10953_ (.I(_04567_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10954_ (.A1(_04890_),
    .A2(_05018_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10955_ (.A1(_02131_),
    .A2(_05037_),
    .B(_05038_),
    .C(_04348_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10956_ (.A1(_00786_),
    .A2(_05018_),
    .B1(_05036_),
    .B2(_05039_),
    .C(_04344_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10957_ (.A1(\as2650.ivec[6] ),
    .A2(_04722_),
    .B1(_04958_),
    .B2(_05018_),
    .C(_04894_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10958_ (.A1(_05015_),
    .A2(_04669_),
    .B1(_05040_),
    .B2(_05041_),
    .C(_04931_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10959_ (.A1(_02238_),
    .A2(_05016_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10960_ (.A1(_04350_),
    .A2(_05042_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10961_ (.I(_05043_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10962_ (.A1(_04370_),
    .A2(_05031_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10963_ (.A1(_04777_),
    .A2(_05043_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10964_ (.A1(_03902_),
    .A2(_05045_),
    .B(_05046_),
    .C(_04699_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(_04387_),
    .A2(_04363_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10966_ (.A1(_02246_),
    .A2(_03992_),
    .B(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10967_ (.A1(_04682_),
    .A2(_05043_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10968_ (.A1(_02571_),
    .A2(_05049_),
    .B(_05050_),
    .C(_03899_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10969_ (.A1(_04615_),
    .A2(_05049_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10970_ (.A1(_04354_),
    .A2(_00880_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10971_ (.A1(_00729_),
    .A2(_05053_),
    .A3(_04768_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10972_ (.A1(_04004_),
    .A2(_05044_),
    .B(_05052_),
    .C(_05054_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10973_ (.A1(_02245_),
    .A2(_05024_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10974_ (.A1(_02245_),
    .A2(_05024_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10975_ (.A1(_05056_),
    .A2(_05057_),
    .B(_00458_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10976_ (.A1(_04619_),
    .A2(_05043_),
    .B(_05058_),
    .C(_04509_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10977_ (.A1(_02589_),
    .A2(_05055_),
    .B(_05059_),
    .C(_00740_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10978_ (.A1(_03711_),
    .A2(_05047_),
    .A3(_05051_),
    .A4(_05060_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10979_ (.A1(_04890_),
    .A2(_05044_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10980_ (.A1(_02155_),
    .A2(_05037_),
    .B(_05062_),
    .C(_03894_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10981_ (.A1(_00786_),
    .A2(_05044_),
    .B1(_05061_),
    .B2(_05063_),
    .C(_04344_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10982_ (.A1(\as2650.ivec[7] ),
    .A2(_04722_),
    .B1(_04958_),
    .B2(_05044_),
    .C(_04609_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10983_ (.A1(_04350_),
    .A2(_04669_),
    .B1(_05064_),
    .B2(_05065_),
    .C(_04931_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10984_ (.I(net69),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10985_ (.A1(net68),
    .A2(_02238_),
    .A3(_05016_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10986_ (.A1(_05066_),
    .A2(_05067_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10987_ (.I(_05068_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10988_ (.A1(_04354_),
    .A2(_05031_),
    .B(_04831_),
    .C(_04355_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10989_ (.A1(_04294_),
    .A2(_05069_),
    .B(_04595_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10990_ (.A1(_02250_),
    .A2(_05057_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10991_ (.A1(_02250_),
    .A2(_05057_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10992_ (.A1(_00456_),
    .A2(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10993_ (.A1(_04823_),
    .A2(_05068_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10994_ (.A1(_05072_),
    .A2(_05074_),
    .B(_05075_),
    .C(_02893_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10995_ (.A1(_02250_),
    .A2(_00551_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10996_ (.A1(_04909_),
    .A2(_05077_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10997_ (.A1(_01024_),
    .A2(_00863_),
    .B1(_03870_),
    .B2(_05068_),
    .C(_05078_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10998_ (.A1(_04497_),
    .A2(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10999_ (.A1(_00739_),
    .A2(_05076_),
    .A3(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11000_ (.A1(_05070_),
    .A2(_05071_),
    .B(_00720_),
    .C(_05081_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11001_ (.A1(_04509_),
    .A2(_05069_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11002_ (.A1(_02580_),
    .A2(_05077_),
    .B(_05083_),
    .C(_00674_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11003_ (.A1(_03711_),
    .A2(_05082_),
    .A3(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11004_ (.A1(_04840_),
    .A2(_05069_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11005_ (.A1(_02176_),
    .A2(_05037_),
    .B(_05085_),
    .C(_05086_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11006_ (.A1(_04611_),
    .A2(_05069_),
    .B1(_05087_),
    .B2(_04564_),
    .C(_04668_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _11007_ (.I(_04666_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11008_ (.A1(_05066_),
    .A2(_04670_),
    .B(_05088_),
    .C(_05089_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11009_ (.I(net90),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11010_ (.A1(_05066_),
    .A2(_05067_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11011_ (.A1(net90),
    .A2(_05091_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11012_ (.I(_05092_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11013_ (.A1(_05090_),
    .A2(_03996_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11014_ (.I0(_05093_),
    .I1(_05094_),
    .S(_03874_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11015_ (.A1(_00456_),
    .A2(_05091_),
    .B(_05074_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11016_ (.A1(net90),
    .A2(_05096_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11017_ (.A1(_04591_),
    .A2(_05092_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11018_ (.A1(_04476_),
    .A2(_00864_),
    .B1(_05094_),
    .B2(_04396_),
    .C(_02586_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11019_ (.A1(_00539_),
    .A2(_05097_),
    .B1(_05098_),
    .B2(_05099_),
    .C(_04595_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11020_ (.A1(_04476_),
    .A2(_04630_),
    .B(_03901_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11021_ (.A1(_04599_),
    .A2(_05093_),
    .B(_00847_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11022_ (.A1(_05101_),
    .A2(_05102_),
    .B(_04331_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11023_ (.A1(_04332_),
    .A2(_05095_),
    .B1(_05100_),
    .B2(_05103_),
    .C(_03987_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11024_ (.A1(_04840_),
    .A2(_05093_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11025_ (.A1(_02193_),
    .A2(_05037_),
    .B(_05104_),
    .C(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11026_ (.A1(_04608_),
    .A2(_05093_),
    .B1(_05106_),
    .B2(_04564_),
    .C(_04668_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11027_ (.A1(_05090_),
    .A2(_04812_),
    .B(_05107_),
    .C(_05089_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11028_ (.A1(_00875_),
    .A2(_03874_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11029_ (.I(_05108_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11030_ (.I(_04124_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11031_ (.A1(_05110_),
    .A2(_01089_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11032_ (.I(_03715_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11033_ (.I(_05112_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11034_ (.A1(_05110_),
    .A2(_01098_),
    .B(_05111_),
    .C(_05113_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11035_ (.I(_04682_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11036_ (.A1(_05115_),
    .A2(_00448_),
    .B(_03894_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11037_ (.A1(net80),
    .A2(_05109_),
    .B(_05114_),
    .C(_05116_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11038_ (.I(_04404_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11039_ (.A1(_02884_),
    .A2(_02881_),
    .B(_05118_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11040_ (.I(_00692_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11041_ (.I(_05120_),
    .Z(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11042_ (.I(_01927_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11043_ (.I(_00930_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11044_ (.A1(_01813_),
    .A2(_05123_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11045_ (.I(_02533_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11046_ (.A1(net88),
    .A2(_05125_),
    .B(_00935_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11047_ (.I(_01926_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11048_ (.A1(_01940_),
    .A2(_04582_),
    .B1(_05124_),
    .B2(_05126_),
    .C(_05127_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11049_ (.I(_02889_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11050_ (.A1(_05122_),
    .A2(_01150_),
    .B(_05128_),
    .C(_05129_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11051_ (.I(_02902_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11052_ (.A1(_05131_),
    .A2(_01110_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11053_ (.A1(_05121_),
    .A2(_05130_),
    .A3(_05132_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11054_ (.I(_02562_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11055_ (.A1(_03841_),
    .A2(_04405_),
    .B1(_05119_),
    .B2(_05133_),
    .C(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11056_ (.A1(_00449_),
    .A2(_04367_),
    .B(_05135_),
    .C(_02922_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11057_ (.A1(_01767_),
    .A2(_01778_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11058_ (.I(_05137_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11059_ (.I(_05138_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11060_ (.A1(\as2650.stack[5][0] ),
    .A2(_03004_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11061_ (.I(_02037_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11062_ (.I(_02035_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11063_ (.A1(\as2650.stack[6][0] ),
    .A2(_05141_),
    .B1(_03088_),
    .B2(\as2650.stack[7][0] ),
    .C1(\as2650.stack[4][0] ),
    .C2(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11064_ (.A1(_05139_),
    .A2(_05140_),
    .A3(_05143_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11065_ (.A1(_02322_),
    .A2(_01772_),
    .B(_02477_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11066_ (.A1(_02202_),
    .A2(_02270_),
    .B(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11067_ (.I(_05146_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11068_ (.I(_05147_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11069_ (.A1(_01799_),
    .A2(_01778_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11070_ (.I(_05149_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11071_ (.I(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11072_ (.A1(\as2650.stack[0][0] ),
    .A2(_02276_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _11073_ (.I(_02091_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11074_ (.A1(\as2650.stack[2][0] ),
    .A2(_05153_),
    .B1(_01805_),
    .B2(\as2650.stack[3][0] ),
    .C1(\as2650.stack[1][0] ),
    .C2(_03331_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11075_ (.A1(_05151_),
    .A2(_05152_),
    .A3(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11076_ (.A1(_05144_),
    .A2(_05148_),
    .A3(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11077_ (.I(_02066_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11078_ (.I(_02165_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11079_ (.A1(\as2650.stack[11][0] ),
    .A2(_05157_),
    .B1(_05158_),
    .B2(\as2650.stack[9][0] ),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11080_ (.I(_02143_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11081_ (.I(_02104_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11082_ (.I(_05137_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11083_ (.A1(\as2650.stack[10][0] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\as2650.stack[8][0] ),
    .C(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11084_ (.A1(_05159_),
    .A2(_05163_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11085_ (.I(_02103_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11086_ (.I(_02077_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11087_ (.A1(\as2650.stack[15][0] ),
    .A2(_05165_),
    .B1(_05166_),
    .B2(\as2650.stack[13][0] ),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11088_ (.I(_02037_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11089_ (.I(_02035_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11090_ (.I(_05149_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11091_ (.A1(\as2650.stack[14][0] ),
    .A2(_05168_),
    .B1(_05169_),
    .B2(\as2650.stack[12][0] ),
    .C(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11092_ (.I(_05147_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11093_ (.A1(_05167_),
    .A2(_05171_),
    .B(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11094_ (.A1(_05164_),
    .A2(_05173_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11095_ (.A1(_05156_),
    .A2(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11096_ (.I(_03757_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11097_ (.A1(_00895_),
    .A2(_00980_),
    .B1(_01025_),
    .B2(_00974_),
    .C(_00591_),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11098_ (.A1(_00982_),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11099_ (.A1(_00564_),
    .A2(_01022_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11100_ (.A1(_04450_),
    .A2(_05179_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11101_ (.A1(_00895_),
    .A2(_00779_),
    .A3(_01022_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11102_ (.A1(_02827_),
    .A2(_03702_),
    .B(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11103_ (.A1(_02792_),
    .A2(_05178_),
    .A3(_05180_),
    .A4(_05182_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11104_ (.A1(_00805_),
    .A2(_02357_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11105_ (.A1(_00840_),
    .A2(_05184_),
    .B(_00895_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11106_ (.A1(_04404_),
    .A2(_04491_),
    .B1(_02524_),
    .B2(_00694_),
    .C(_00839_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(_00580_),
    .A2(_03713_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11108_ (.A1(_00783_),
    .A2(_05183_),
    .B1(_05185_),
    .B2(_05186_),
    .C(_05187_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11109_ (.A1(_02811_),
    .A2(_00688_),
    .A3(_00956_),
    .A4(_02537_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11110_ (.A1(_02798_),
    .A2(_02800_),
    .A3(_02803_),
    .A4(_03124_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11111_ (.A1(_02811_),
    .A2(_00509_),
    .A3(_00625_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11112_ (.A1(_02859_),
    .A2(_00530_),
    .A3(_00632_),
    .A4(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11113_ (.A1(_00819_),
    .A2(_05189_),
    .B(_05190_),
    .C(_05192_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11114_ (.A1(_05176_),
    .A2(_05188_),
    .B(_05193_),
    .C(_02789_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11115_ (.I(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11116_ (.I(_05195_),
    .Z(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11117_ (.A1(_05117_),
    .A2(_05136_),
    .B1(_05175_),
    .B2(_04481_),
    .C(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11118_ (.I(_05194_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11119_ (.I(_05198_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11120_ (.I(_02998_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11121_ (.A1(_01139_),
    .A2(_05199_),
    .B(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11122_ (.A1(_05197_),
    .A2(_05201_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11123_ (.I(_05176_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11124_ (.A1(_04168_),
    .A2(_01229_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11125_ (.A1(_04028_),
    .A2(_01200_),
    .B(_00907_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11126_ (.A1(_04508_),
    .A2(_02884_),
    .B1(_05203_),
    .B2(_05204_),
    .C(_03893_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11127_ (.A1(_01188_),
    .A2(_05108_),
    .B(_05205_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11128_ (.A1(_01830_),
    .A2(_00930_),
    .B(_02572_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11129_ (.A1(_02322_),
    .A2(_00931_),
    .B(_05207_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11130_ (.A1(_01939_),
    .A2(_04661_),
    .B(_05208_),
    .C(_01927_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11131_ (.A1(_05127_),
    .A2(_01237_),
    .B(_05209_),
    .C(_02889_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11132_ (.A1(_00787_),
    .A2(_05809_),
    .B(_05120_),
    .C(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11133_ (.A1(_01267_),
    .A2(_05121_),
    .B(_05211_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11134_ (.A1(_02905_),
    .A2(_05212_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11135_ (.A1(_04537_),
    .A2(_02861_),
    .B(_05010_),
    .C(_05213_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11136_ (.A1(_00451_),
    .A2(_00464_),
    .B(_05206_),
    .C(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11137_ (.I(_05147_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11138_ (.I(_02034_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11139_ (.I(_02112_),
    .Z(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11140_ (.A1(\as2650.stack[7][1] ),
    .A2(_05217_),
    .B1(_05218_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11141_ (.A1(\as2650.stack[6][1] ),
    .A2(_05153_),
    .B1(_02375_),
    .B2(\as2650.stack[4][1] ),
    .C(_05150_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11142_ (.A1(_05219_),
    .A2(_05220_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11143_ (.I(_05149_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(\as2650.stack[1][1] ),
    .A2(_05166_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11145_ (.I(_01993_),
    .Z(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11146_ (.I(_02127_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11147_ (.I(_02023_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11148_ (.A1(\as2650.stack[2][1] ),
    .A2(_05224_),
    .B1(_05225_),
    .B2(\as2650.stack[3][1] ),
    .C1(\as2650.stack[0][1] ),
    .C2(_05226_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11149_ (.A1(_05222_),
    .A2(_05223_),
    .A3(_05227_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(_05221_),
    .A2(_05228_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11151_ (.I(_05137_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(\as2650.stack[13][1] ),
    .A2(_05218_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11153_ (.I(_02083_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11154_ (.I(_01982_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11155_ (.A1(\as2650.stack[14][1] ),
    .A2(_05224_),
    .B1(_05232_),
    .B2(\as2650.stack[15][1] ),
    .C1(\as2650.stack[12][1] ),
    .C2(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11156_ (.A1(_05230_),
    .A2(_05231_),
    .A3(_05234_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11157_ (.A1(\as2650.stack[9][1] ),
    .A2(_03331_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11158_ (.A1(\as2650.stack[10][1] ),
    .A2(_02079_),
    .B1(_05232_),
    .B2(\as2650.stack[11][1] ),
    .C1(\as2650.stack[8][1] ),
    .C2(_05233_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11159_ (.A1(_05222_),
    .A2(_05236_),
    .A3(_05237_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11160_ (.I(_05147_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11161_ (.A1(_05235_),
    .A2(_05238_),
    .B(_05239_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11162_ (.I(_05176_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11163_ (.A1(_05216_),
    .A2(_05229_),
    .B(_05240_),
    .C(_05241_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11164_ (.A1(_05202_),
    .A2(_05215_),
    .B(_05242_),
    .C(_05196_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11165_ (.A1(_02676_),
    .A2(_05199_),
    .B(_05200_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11166_ (.A1(_05243_),
    .A2(_05244_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11167_ (.I(_00579_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11168_ (.A1(_05245_),
    .A2(_01275_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11169_ (.A1(_05110_),
    .A2(_01269_),
    .B(_05112_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11170_ (.A1(_04406_),
    .A2(_01267_),
    .B(_03893_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11171_ (.A1(_01299_),
    .A2(_05108_),
    .B1(_05246_),
    .B2(_05247_),
    .C(_05248_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11172_ (.I(_02860_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11173_ (.A1(_01772_),
    .A2(_03758_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11174_ (.A1(_01844_),
    .A2(_05125_),
    .B(_01939_),
    .C(_05251_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11175_ (.A1(_00935_),
    .A2(_04719_),
    .B(_05252_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11176_ (.A1(_02892_),
    .A2(_05127_),
    .A3(_05253_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11177_ (.A1(_01927_),
    .A2(_01313_),
    .B(_00692_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11178_ (.A1(_01249_),
    .A2(_02902_),
    .B(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11179_ (.A1(_01404_),
    .A2(_02880_),
    .B1(_05254_),
    .B2(_05256_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11180_ (.A1(_02905_),
    .A2(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11181_ (.A1(_02868_),
    .A2(_05250_),
    .B(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11182_ (.A1(_00443_),
    .A2(_03922_),
    .B1(_05010_),
    .B2(_05259_),
    .C(_04480_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11183_ (.A1(\as2650.stack[7][2] ),
    .A2(_03088_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11184_ (.I(_02151_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11185_ (.A1(\as2650.stack[5][2] ),
    .A2(_05262_),
    .B1(_05233_),
    .B2(\as2650.stack[4][2] ),
    .C1(\as2650.stack[6][2] ),
    .C2(_05224_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11186_ (.A1(_05230_),
    .A2(_05261_),
    .A3(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(\as2650.stack[2][2] ),
    .A2(_05141_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11188_ (.A1(\as2650.stack[1][2] ),
    .A2(_05262_),
    .B1(_02085_),
    .B2(\as2650.stack[0][2] ),
    .C1(\as2650.stack[3][2] ),
    .C2(_05232_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11189_ (.A1(_05222_),
    .A2(_05265_),
    .A3(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11190_ (.A1(_05264_),
    .A2(_05267_),
    .ZN(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11191_ (.A1(\as2650.stack[12][2] ),
    .A2(_02375_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11192_ (.A1(\as2650.stack[14][2] ),
    .A2(_02079_),
    .B1(_02084_),
    .B2(\as2650.stack[15][2] ),
    .C1(\as2650.stack[13][2] ),
    .C2(_02087_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11193_ (.A1(_05162_),
    .A2(_05269_),
    .A3(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11194_ (.I(_01962_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11195_ (.A1(\as2650.stack[8][2] ),
    .A2(_05272_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11196_ (.A1(\as2650.stack[10][2] ),
    .A2(_02169_),
    .B1(_02119_),
    .B2(\as2650.stack[11][2] ),
    .C1(\as2650.stack[9][2] ),
    .C2(_02087_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11197_ (.A1(_05170_),
    .A2(_05273_),
    .A3(_05274_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11198_ (.A1(_05271_),
    .A2(_05275_),
    .B(_05172_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11199_ (.A1(_05148_),
    .A2(_05268_),
    .B(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11200_ (.I(_05195_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11201_ (.A1(_05249_),
    .A2(_05260_),
    .B1(_05277_),
    .B2(_02933_),
    .C(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11202_ (.A1(_01847_),
    .A2(_05196_),
    .B(_05279_),
    .C(_05089_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11203_ (.A1(_04124_),
    .A2(_01362_),
    .B(_05112_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11204_ (.A1(_04063_),
    .A2(_03206_),
    .B(_05280_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11205_ (.A1(_04406_),
    .A2(_01404_),
    .B(_05281_),
    .C(_00785_),
    .ZN(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11206_ (.A1(_02844_),
    .A2(_05108_),
    .B(_05282_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11207_ (.I(_05120_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11208_ (.A1(_01780_),
    .A2(_05125_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11209_ (.A1(_01107_),
    .A2(_05123_),
    .B(_02572_),
    .ZN(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11210_ (.A1(_05285_),
    .A2(_05286_),
    .B(_02902_),
    .C(_00957_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11211_ (.A1(_00936_),
    .A2(_04741_),
    .B(_05287_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11212_ (.A1(_01267_),
    .A2(_05131_),
    .B1(_00957_),
    .B2(_01385_),
    .C(_02880_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11213_ (.A1(_05288_),
    .A2(_05289_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11214_ (.A1(_02883_),
    .A2(_05284_),
    .B(_05290_),
    .C(_05250_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11215_ (.I(_02872_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11216_ (.A1(_05292_),
    .A2(_05118_),
    .B(_02562_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11217_ (.A1(_00428_),
    .A2(_00463_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11218_ (.A1(_05291_),
    .A2(_05293_),
    .B(_04480_),
    .C(_05294_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(\as2650.stack[6][3] ),
    .A2(_05141_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11220_ (.A1(\as2650.stack[5][3] ),
    .A2(_05262_),
    .B1(_05233_),
    .B2(\as2650.stack[4][3] ),
    .C1(\as2650.stack[7][3] ),
    .C2(_05232_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11221_ (.A1(_05162_),
    .A2(_05296_),
    .A3(_05297_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11222_ (.I(_01804_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11223_ (.I(_01986_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11224_ (.A1(\as2650.stack[3][3] ),
    .A2(_05299_),
    .B1(_05300_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11225_ (.A1(\as2650.stack[2][3] ),
    .A2(_05224_),
    .B1(_05226_),
    .B2(\as2650.stack[0][3] ),
    .C(_05138_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11226_ (.A1(_05301_),
    .A2(_05302_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11227_ (.A1(_05298_),
    .A2(_05303_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11228_ (.A1(\as2650.stack[10][3] ),
    .A2(_05153_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11229_ (.A1(\as2650.stack[9][3] ),
    .A2(_02087_),
    .B1(_02085_),
    .B2(\as2650.stack[8][3] ),
    .C1(\as2650.stack[11][3] ),
    .C2(_02084_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11230_ (.A1(_05222_),
    .A2(_05305_),
    .A3(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11231_ (.I(_02091_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11232_ (.A1(\as2650.stack[14][3] ),
    .A2(_05308_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11233_ (.A1(\as2650.stack[13][3] ),
    .A2(_02122_),
    .B1(_02085_),
    .B2(\as2650.stack[12][3] ),
    .C1(\as2650.stack[15][3] ),
    .C2(_02084_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11234_ (.A1(_05162_),
    .A2(_05309_),
    .A3(_05310_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11235_ (.A1(_05307_),
    .A2(_05311_),
    .B(_05172_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11236_ (.A1(_05148_),
    .A2(_05304_),
    .B(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11237_ (.I(_00798_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11238_ (.A1(_05283_),
    .A2(_05295_),
    .B1(_05313_),
    .B2(_05314_),
    .C(_05195_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11239_ (.A1(_01354_),
    .A2(_05196_),
    .B(_05315_),
    .C(_05089_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11240_ (.A1(_03969_),
    .A2(_03223_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11241_ (.A1(_05245_),
    .A2(_01428_),
    .B(_05316_),
    .C(_05113_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11242_ (.A1(_05115_),
    .A2(_02883_),
    .B(_03894_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11243_ (.A1(_01456_),
    .A2(_05109_),
    .B(_05317_),
    .C(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11244_ (.A1(_05122_),
    .A2(_01634_),
    .B(_05129_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11245_ (.I(net74),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11246_ (.A1(_05321_),
    .A2(_00932_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11247_ (.A1(_03233_),
    .A2(_00932_),
    .B(_02530_),
    .C(_05322_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11248_ (.A1(_02574_),
    .A2(_04809_),
    .B(_05320_),
    .C(_05323_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11249_ (.A1(_03187_),
    .A2(_02957_),
    .B(_05121_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11250_ (.A1(_01570_),
    .A2(_05284_),
    .B1(_05324_),
    .B2(_05325_),
    .C(_05250_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11251_ (.A1(_02876_),
    .A2(_04405_),
    .B(_05134_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11252_ (.A1(_00432_),
    .A2(_03922_),
    .B1(_05326_),
    .B2(_05327_),
    .C(_02922_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11253_ (.A1(\as2650.stack[4][4] ),
    .A2(_02276_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11254_ (.A1(\as2650.stack[6][4] ),
    .A2(_05153_),
    .B1(_01805_),
    .B2(\as2650.stack[7][4] ),
    .C1(\as2650.stack[5][4] ),
    .C2(_05300_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11255_ (.A1(_05139_),
    .A2(_05329_),
    .A3(_05330_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11256_ (.A1(\as2650.stack[2][4] ),
    .A2(_05160_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11257_ (.A1(\as2650.stack[1][4] ),
    .A2(_05300_),
    .B1(_05142_),
    .B2(\as2650.stack[0][4] ),
    .C1(\as2650.stack[3][4] ),
    .C2(_01805_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11258_ (.A1(_05151_),
    .A2(_05332_),
    .A3(_05333_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11259_ (.A1(_05148_),
    .A2(_05331_),
    .A3(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11260_ (.A1(\as2650.stack[11][4] ),
    .A2(_05157_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11261_ (.A1(\as2650.stack[9][4] ),
    .A2(_05218_),
    .B1(_05142_),
    .B2(\as2650.stack[8][4] ),
    .C1(\as2650.stack[10][4] ),
    .C2(_05141_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11262_ (.A1(_05151_),
    .A2(_05336_),
    .A3(_05337_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11263_ (.A1(\as2650.stack[15][4] ),
    .A2(_05165_),
    .B1(_05166_),
    .B2(\as2650.stack[13][4] ),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11264_ (.A1(\as2650.stack[14][4] ),
    .A2(_05168_),
    .B1(_05142_),
    .B2(\as2650.stack[12][4] ),
    .C(_05150_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11265_ (.A1(_05339_),
    .A2(_05340_),
    .B(_05172_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11266_ (.A1(_05338_),
    .A2(_05341_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11267_ (.A1(_05335_),
    .A2(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11268_ (.A1(_05319_),
    .A2(_05328_),
    .B1(_05343_),
    .B2(_04481_),
    .C(_05278_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11269_ (.A1(_03647_),
    .A2(_05199_),
    .B(_05200_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11270_ (.A1(_05344_),
    .A2(_05345_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11271_ (.A1(_05110_),
    .A2(_01509_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11272_ (.A1(_05245_),
    .A2(_01493_),
    .B(_05113_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11273_ (.A1(_05115_),
    .A2(_01570_),
    .B(_03719_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11274_ (.A1(_01534_),
    .A2(_05109_),
    .B1(_05346_),
    .B2(_05347_),
    .C(_05348_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11275_ (.A1(_02573_),
    .A2(_04857_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(_01888_),
    .A2(_00931_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11277_ (.A1(_02593_),
    .A2(_05123_),
    .B(_01940_),
    .C(_05351_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11278_ (.A1(_01928_),
    .A2(_05350_),
    .A3(_05352_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11279_ (.A1(_05122_),
    .A2(_01631_),
    .B(_05353_),
    .C(_00626_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11280_ (.A1(_01670_),
    .A2(_02881_),
    .B1(_05131_),
    .B2(_02883_),
    .C(_04404_),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11281_ (.A1(_02584_),
    .A2(_05118_),
    .B1(_05354_),
    .B2(_05355_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11282_ (.I(_05176_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11283_ (.A1(_05134_),
    .A2(_05356_),
    .B(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11284_ (.A1(_00425_),
    .A2(_04367_),
    .B(_05358_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11285_ (.A1(\as2650.stack[7][5] ),
    .A2(_05217_),
    .B1(_05166_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11286_ (.A1(\as2650.stack[6][5] ),
    .A2(_05168_),
    .B1(_05169_),
    .B2(\as2650.stack[4][5] ),
    .C(_05170_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(_05360_),
    .A2(_05361_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11288_ (.I(_05150_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11289_ (.A1(\as2650.stack[1][5] ),
    .A2(_05158_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11290_ (.A1(\as2650.stack[2][5] ),
    .A2(_05308_),
    .B1(_05299_),
    .B2(\as2650.stack[3][5] ),
    .C1(\as2650.stack[0][5] ),
    .C2(_05272_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11291_ (.A1(_05363_),
    .A2(_05364_),
    .A3(_05365_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11292_ (.A1(_05362_),
    .A2(_05366_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11293_ (.A1(\as2650.stack[10][5] ),
    .A2(_05160_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11294_ (.I(_02151_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11295_ (.A1(\as2650.stack[9][5] ),
    .A2(_05369_),
    .B1(_05272_),
    .B2(\as2650.stack[8][5] ),
    .C1(\as2650.stack[11][5] ),
    .C2(_05299_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11296_ (.A1(_05363_),
    .A2(_05368_),
    .A3(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11297_ (.I(_02143_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11298_ (.A1(\as2650.stack[14][5] ),
    .A2(_05372_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11299_ (.A1(\as2650.stack[13][5] ),
    .A2(_05369_),
    .B1(_05226_),
    .B2(\as2650.stack[12][5] ),
    .C1(\as2650.stack[15][5] ),
    .C2(_05225_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11300_ (.A1(_05230_),
    .A2(_05373_),
    .A3(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11301_ (.A1(_05371_),
    .A2(_05375_),
    .B(_05239_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11302_ (.A1(_05216_),
    .A2(_05367_),
    .B(_05376_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11303_ (.A1(_05349_),
    .A2(_05359_),
    .B1(_05377_),
    .B2(_04481_),
    .C(_05278_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11304_ (.A1(_03316_),
    .A2(_05198_),
    .B(_05200_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11305_ (.A1(_05378_),
    .A2(_05379_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11306_ (.A1(_03969_),
    .A2(_01592_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11307_ (.A1(_05245_),
    .A2(_01597_),
    .B(_05380_),
    .C(_05113_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11308_ (.A1(_05115_),
    .A2(_01670_),
    .B(_03719_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11309_ (.A1(_01622_),
    .A2(_05109_),
    .B(_05381_),
    .C(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(net29),
    .A2(_05125_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11311_ (.A1(_02897_),
    .A2(_00932_),
    .B(_02530_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11312_ (.A1(_01928_),
    .A2(_02256_),
    .B(_05120_),
    .C(_02892_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11313_ (.A1(_02574_),
    .A2(_02921_),
    .B1(_05384_),
    .B2(_05385_),
    .C(_05386_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11314_ (.I(_01579_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11315_ (.A1(_05388_),
    .A2(_05121_),
    .B1(_05129_),
    .B2(_01413_),
    .C(_02905_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11316_ (.A1(_04524_),
    .A2(_05250_),
    .B1(_05387_),
    .B2(_05389_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11317_ (.A1(_00422_),
    .A2(_03922_),
    .B1(_05010_),
    .B2(_05390_),
    .C(_02922_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11318_ (.A1(\as2650.stack[7][6] ),
    .A2(_05165_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11319_ (.A1(\as2650.stack[5][6] ),
    .A2(_05369_),
    .B1(_02375_),
    .B2(\as2650.stack[4][6] ),
    .C1(\as2650.stack[6][6] ),
    .C2(_05308_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11320_ (.A1(_05139_),
    .A2(_05392_),
    .A3(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11321_ (.A1(\as2650.stack[0][6] ),
    .A2(_05161_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11322_ (.A1(\as2650.stack[2][6] ),
    .A2(_05308_),
    .B1(_05299_),
    .B2(\as2650.stack[3][6] ),
    .C1(\as2650.stack[1][6] ),
    .C2(_05300_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11323_ (.A1(_05363_),
    .A2(_05395_),
    .A3(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11324_ (.A1(_05394_),
    .A2(_05397_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11325_ (.A1(\as2650.stack[10][6] ),
    .A2(_05372_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11326_ (.A1(\as2650.stack[9][6] ),
    .A2(_05369_),
    .B1(_05272_),
    .B2(\as2650.stack[8][6] ),
    .C1(\as2650.stack[11][6] ),
    .C2(_05225_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11327_ (.A1(_05363_),
    .A2(_05399_),
    .A3(_05400_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11328_ (.A1(\as2650.stack[14][6] ),
    .A2(_05168_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11329_ (.A1(\as2650.stack[13][6] ),
    .A2(_05262_),
    .B1(_05226_),
    .B2(\as2650.stack[12][6] ),
    .C1(\as2650.stack[15][6] ),
    .C2(_05225_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11330_ (.A1(_05230_),
    .A2(_05402_),
    .A3(_05403_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11331_ (.A1(_05401_),
    .A2(_05404_),
    .B(_05239_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11332_ (.A1(_05216_),
    .A2(_05398_),
    .B(_05405_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11333_ (.A1(_05383_),
    .A2(_05391_),
    .B1(_05406_),
    .B2(_02933_),
    .C(_05278_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11334_ (.I(_02998_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11335_ (.A1(_03672_),
    .A2(_05198_),
    .B(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11336_ (.A1(_05407_),
    .A2(_05409_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11337_ (.A1(_00778_),
    .A2(_02581_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11338_ (.A1(_04063_),
    .A2(_01692_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11339_ (.A1(_04028_),
    .A2(_01687_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11340_ (.A1(_05112_),
    .A2(_05411_),
    .A3(_05412_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11341_ (.A1(_00571_),
    .A2(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11342_ (.A1(_02854_),
    .A2(_05388_),
    .B1(_02928_),
    .B2(_05410_),
    .C(_05414_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11343_ (.A1(_02573_),
    .A2(_02956_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11344_ (.A1(_05717_),
    .A2(_00931_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11345_ (.A1(net77),
    .A2(_05123_),
    .B(_00935_),
    .C(_05417_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11346_ (.A1(_05127_),
    .A2(_05416_),
    .A3(_05418_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11347_ (.A1(_05122_),
    .A2(_03462_),
    .B(_05419_),
    .C(_05129_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11348_ (.A1(_02881_),
    .A2(_01673_),
    .B1(_02903_),
    .B2(_05420_),
    .C(_05118_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11349_ (.A1(_00554_),
    .A2(_04405_),
    .B(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11350_ (.A1(_05840_),
    .A2(_00464_),
    .B1(_05134_),
    .B2(_05422_),
    .C(_05241_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11351_ (.A1(\as2650.stack[13][7] ),
    .A2(_03004_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11352_ (.A1(\as2650.stack[14][7] ),
    .A2(_05372_),
    .B1(_05217_),
    .B2(\as2650.stack[15][7] ),
    .C1(\as2650.stack[12][7] ),
    .C2(_05169_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11353_ (.A1(_05139_),
    .A2(_05424_),
    .A3(_05425_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11354_ (.A1(\as2650.stack[11][7] ),
    .A2(_05165_),
    .B1(_05158_),
    .B2(\as2650.stack[9][7] ),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11355_ (.A1(\as2650.stack[10][7] ),
    .A2(_05372_),
    .B1(_05161_),
    .B2(\as2650.stack[8][7] ),
    .C(_05138_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11356_ (.A1(_05427_),
    .A2(_05428_),
    .B(_05239_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11357_ (.A1(_05426_),
    .A2(_05429_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11358_ (.A1(\as2650.stack[7][7] ),
    .A2(_05157_),
    .B1(_05158_),
    .B2(\as2650.stack[5][7] ),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11359_ (.A1(\as2650.stack[6][7] ),
    .A2(_05160_),
    .B1(_05161_),
    .B2(\as2650.stack[4][7] ),
    .C(_05170_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11360_ (.A1(_05431_),
    .A2(_05432_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11361_ (.A1(\as2650.stack[2][7] ),
    .A2(_02424_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11362_ (.A1(\as2650.stack[1][7] ),
    .A2(_05218_),
    .B1(_05169_),
    .B2(\as2650.stack[0][7] ),
    .C1(\as2650.stack[3][7] ),
    .C2(_05217_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11363_ (.A1(_05151_),
    .A2(_05434_),
    .A3(_05435_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11364_ (.A1(_05216_),
    .A2(_05433_),
    .A3(_05436_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11365_ (.A1(_05314_),
    .A2(_05430_),
    .A3(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11366_ (.A1(_05415_),
    .A2(_05423_),
    .B(_05438_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11367_ (.A1(_01678_),
    .A2(_05198_),
    .B(_04381_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11368_ (.A1(_05199_),
    .A2(_05439_),
    .B(_05440_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11369_ (.A1(_01932_),
    .A2(_02360_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11370_ (.A1(_01100_),
    .A2(_04497_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11371_ (.A1(_00922_),
    .A2(_05442_),
    .B1(_04941_),
    .B2(_02203_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11372_ (.A1(_05441_),
    .A2(_04498_),
    .B(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11373_ (.A1(_04566_),
    .A2(_05444_),
    .B(_05202_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11374_ (.A1(_00933_),
    .A2(_02777_),
    .B(_02598_),
    .ZN(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11375_ (.A1(_04416_),
    .A2(_04418_),
    .B(_04421_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11376_ (.A1(_00765_),
    .A2(_00599_),
    .A3(_04422_),
    .A4(_04461_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11377_ (.I(_02780_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11378_ (.A1(_00839_),
    .A2(_02566_),
    .B(_05449_),
    .C(_00735_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11379_ (.A1(_00537_),
    .A2(_00769_),
    .B(_05450_),
    .C(_00718_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11380_ (.A1(_00986_),
    .A2(_04420_),
    .A3(_03731_),
    .A4(_04448_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11381_ (.A1(_02559_),
    .A2(_05451_),
    .B(_05452_),
    .C(_04426_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11382_ (.A1(_00471_),
    .A2(_05824_),
    .B(_00516_),
    .C(_00789_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11383_ (.A1(_04556_),
    .A2(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11384_ (.A1(_00520_),
    .A2(_05455_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11385_ (.A1(_02556_),
    .A2(_05453_),
    .A3(_05456_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11386_ (.A1(_02561_),
    .A2(_05448_),
    .A3(_05457_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11387_ (.A1(_02528_),
    .A2(_02551_),
    .A3(_05447_),
    .A4(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11388_ (.I(_05459_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11389_ (.A1(_05445_),
    .A2(_05446_),
    .B(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11390_ (.A1(_04840_),
    .A2(_05444_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11391_ (.A1(_05241_),
    .A2(_05462_),
    .B(_02597_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11392_ (.A1(_05460_),
    .A2(_05463_),
    .B(_02203_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11393_ (.A1(_04060_),
    .A2(_05464_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11394_ (.A1(_01813_),
    .A2(_05461_),
    .B(_05465_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11395_ (.I(\as2650.r123_2[3][0] ),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11396_ (.I(_05466_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11397_ (.I(\as2650.r123_2[3][1] ),
    .Z(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11398_ (.I(_05467_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11399_ (.I(\as2650.r123_2[3][2] ),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11400_ (.I(_05468_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11401_ (.I(\as2650.r123_2[3][3] ),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11402_ (.I(_05469_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11403_ (.I(\as2650.r123_2[3][4] ),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11404_ (.I(_05470_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11405_ (.I(\as2650.r123_2[3][5] ),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11406_ (.I(_05471_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11407_ (.I(\as2650.r123_2[3][6] ),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11408_ (.I(_05472_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11409_ (.I(\as2650.r123_2[3][7] ),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11410_ (.I(_05473_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11411_ (.A1(_02628_),
    .A2(_01815_),
    .A3(_02271_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11412_ (.I(_05474_),
    .Z(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11413_ (.I(_05475_),
    .Z(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11414_ (.A1(\as2650.stack[9][8] ),
    .A2(_05475_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11415_ (.A1(_01765_),
    .A2(_01948_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11416_ (.I(_05478_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11417_ (.I(_05479_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11418_ (.A1(_02718_),
    .A2(_05476_),
    .B(_05477_),
    .C(_05480_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11419_ (.I(_05474_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11420_ (.A1(\as2650.stack[9][9] ),
    .A2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11421_ (.A1(_02726_),
    .A2(_05476_),
    .B(_05480_),
    .C(_05482_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11422_ (.I(_05474_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11423_ (.A1(\as2650.stack[9][10] ),
    .A2(_05483_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11424_ (.A1(_02729_),
    .A2(_05476_),
    .B(_05480_),
    .C(_05484_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11425_ (.A1(\as2650.stack[9][11] ),
    .A2(_05483_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11426_ (.A1(_02732_),
    .A2(_05476_),
    .B(_05480_),
    .C(_05485_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11427_ (.I(_05475_),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11428_ (.I(_05479_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11429_ (.A1(\as2650.stack[9][12] ),
    .A2(_05483_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11430_ (.A1(_02734_),
    .A2(_05486_),
    .B(_05487_),
    .C(_05488_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11431_ (.A1(\as2650.stack[9][13] ),
    .A2(_05483_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11432_ (.A1(_02738_),
    .A2(_05486_),
    .B(_05487_),
    .C(_05489_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11433_ (.A1(\as2650.stack[9][14] ),
    .A2(_05475_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11434_ (.A1(_02740_),
    .A2(_05486_),
    .B(_05487_),
    .C(_05490_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11435_ (.I(_05478_),
    .Z(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11436_ (.I(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11437_ (.A1(_02275_),
    .A2(_05157_),
    .A3(_02277_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11438_ (.I(_05493_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11439_ (.A1(\as2650.stack[9][0] ),
    .A2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11440_ (.I(_05474_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11441_ (.A1(_01825_),
    .A2(_05496_),
    .B(_05487_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11442_ (.A1(_03575_),
    .A2(_05492_),
    .B1(_05495_),
    .B2(_05497_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11443_ (.A1(_03037_),
    .A2(_05486_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11444_ (.I(_05493_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11445_ (.I(_05479_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11446_ (.A1(\as2650.stack[9][1] ),
    .A2(_05499_),
    .B(_05500_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11447_ (.A1(_01831_),
    .A2(_05492_),
    .B1(_05498_),
    .B2(_05501_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11448_ (.A1(\as2650.stack[9][2] ),
    .A2(_05494_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11449_ (.A1(_01858_),
    .A2(_05481_),
    .B(_05500_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11450_ (.A1(_01845_),
    .A2(_05492_),
    .B1(_05502_),
    .B2(_05503_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11451_ (.A1(_03100_),
    .A2(_05496_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11452_ (.A1(\as2650.stack[9][3] ),
    .A2(_05499_),
    .B(_05500_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11453_ (.A1(_03589_),
    .A2(_05492_),
    .B1(_05504_),
    .B2(_05505_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11454_ (.I(_05479_),
    .Z(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11455_ (.A1(_01884_),
    .A2(_05496_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11456_ (.A1(\as2650.stack[9][4] ),
    .A2(_05499_),
    .B(_05500_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11457_ (.A1(_01873_),
    .A2(_05506_),
    .B1(_05507_),
    .B2(_05508_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11458_ (.A1(\as2650.stack[9][5] ),
    .A2(_05494_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11459_ (.A1(_01899_),
    .A2(_05481_),
    .B(_05491_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11460_ (.A1(_01889_),
    .A2(_05506_),
    .B1(_05509_),
    .B2(_05510_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11461_ (.A1(\as2650.stack[9][6] ),
    .A2(_05494_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11462_ (.A1(_03354_),
    .A2(_05481_),
    .B(_05491_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11463_ (.A1(_01902_),
    .A2(_05506_),
    .B1(_05511_),
    .B2(_05512_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11464_ (.A1(_02314_),
    .A2(_05496_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11465_ (.A1(\as2650.stack[9][7] ),
    .A2(_05499_),
    .B(_05491_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11466_ (.A1(_03599_),
    .A2(_05506_),
    .B1(_05513_),
    .B2(_05514_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11467_ (.A1(_00479_),
    .A2(_01029_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11468_ (.I(_05515_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11469_ (.I(_05516_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11470_ (.A1(_01153_),
    .A2(_05515_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11471_ (.I(_05518_),
    .Z(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11472_ (.A1(\as2650.r123[2][0] ),
    .A2(_05519_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11473_ (.I(_01144_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11474_ (.A1(_05521_),
    .A2(_03401_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11475_ (.A1(_01136_),
    .A2(_05517_),
    .B(_05520_),
    .C(_05522_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11476_ (.A1(_05521_),
    .A2(_03438_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11477_ (.I(_05518_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11478_ (.A1(\as2650.r123[2][1] ),
    .A2(_05524_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11479_ (.A1(_01232_),
    .A2(_05517_),
    .B(_05523_),
    .C(_05525_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11480_ (.A1(_05521_),
    .A2(_03477_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11481_ (.A1(\as2650.r123[2][2] ),
    .A2(_05524_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11482_ (.A1(_01301_),
    .A2(_05517_),
    .B(_05526_),
    .C(_05527_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11483_ (.A1(_05521_),
    .A2(_03506_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11484_ (.A1(\as2650.r123[2][3] ),
    .A2(_05524_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11485_ (.A1(_01370_),
    .A2(_05517_),
    .B(_05528_),
    .C(_05529_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11486_ (.I(_05515_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11487_ (.A1(_01457_),
    .A2(_05530_),
    .B1(_05519_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11488_ (.A1(_01461_),
    .A2(_03521_),
    .B(_05531_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11489_ (.A1(_01244_),
    .A2(_03534_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11490_ (.A1(\as2650.r123[2][5] ),
    .A2(_05524_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11491_ (.A1(_01536_),
    .A2(_05516_),
    .B(_05532_),
    .C(_05533_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(_01244_),
    .A2(_03543_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11493_ (.A1(\as2650.r123[2][6] ),
    .A2(_05519_),
    .ZN(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11494_ (.A1(_01624_),
    .A2(_05516_),
    .B(_05534_),
    .C(_05535_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11495_ (.A1(_03546_),
    .A2(_03547_),
    .A3(_03548_),
    .B(_01144_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11496_ (.A1(\as2650.r123[2][7] ),
    .A2(_05519_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11497_ (.A1(_01718_),
    .A2(_05516_),
    .B(_05536_),
    .C(_05537_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11498_ (.A1(_00623_),
    .A2(_04450_),
    .A3(_05179_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11499_ (.A1(_00572_),
    .A2(_00574_),
    .B(_00577_),
    .C(_00580_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11500_ (.A1(_04388_),
    .A2(_05539_),
    .B(_03714_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11501_ (.A1(_00790_),
    .A2(_02852_),
    .A3(_03709_),
    .B(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11502_ (.A1(_03787_),
    .A2(_05538_),
    .B(_05541_),
    .C(_03705_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11503_ (.I(_05542_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11504_ (.A1(_00784_),
    .A2(_01025_),
    .Z(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11505_ (.I(_05544_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11506_ (.I(_05544_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11507_ (.A1(_01217_),
    .A2(_05546_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11508_ (.A1(_01138_),
    .A2(_05545_),
    .B(_05547_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11509_ (.I(_05542_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11510_ (.A1(net43),
    .A2(_05549_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11511_ (.I(_04666_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11512_ (.A1(_05543_),
    .A2(_05548_),
    .B(_05550_),
    .C(_05551_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11513_ (.A1(_02884_),
    .A2(_05546_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11514_ (.A1(_02676_),
    .A2(_05545_),
    .B(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11515_ (.A1(net44),
    .A2(_05549_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11516_ (.A1(_05543_),
    .A2(_05553_),
    .B(_05554_),
    .C(_05551_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11517_ (.A1(_01345_),
    .A2(_05546_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11518_ (.A1(_01247_),
    .A2(_05545_),
    .B(_05555_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11519_ (.A1(net45),
    .A2(_05549_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11520_ (.A1(_05543_),
    .A2(_05556_),
    .B(_05557_),
    .C(_05551_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11521_ (.A1(_03187_),
    .A2(_05546_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11522_ (.A1(_02133_),
    .A2(_05545_),
    .B(_05558_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11523_ (.A1(net46),
    .A2(_05549_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11524_ (.A1(_05543_),
    .A2(_05559_),
    .B(_05560_),
    .C(_05551_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11525_ (.I(_05542_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11526_ (.I(_05544_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_05544_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11528_ (.A1(_01497_),
    .A2(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11529_ (.A1(_03647_),
    .A2(_05562_),
    .B(_05564_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11530_ (.I(_05542_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11531_ (.A1(net47),
    .A2(_05566_),
    .ZN(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11532_ (.I(_04666_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11533_ (.A1(_05561_),
    .A2(_05565_),
    .B(_05567_),
    .C(_05568_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11534_ (.A1(_01413_),
    .A2(_05563_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11535_ (.A1(_03316_),
    .A2(_05562_),
    .B(_05569_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11536_ (.A1(net21),
    .A2(_05566_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11537_ (.A1(_05561_),
    .A2(_05570_),
    .B(_05571_),
    .C(_05568_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11538_ (.A1(_02886_),
    .A2(_05563_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11539_ (.A1(_03672_),
    .A2(_05562_),
    .B(_05572_),
    .ZN(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11540_ (.A1(net22),
    .A2(_05566_),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11541_ (.A1(_05561_),
    .A2(_05573_),
    .B(_05574_),
    .C(_05568_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11542_ (.A1(_05388_),
    .A2(_05563_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11543_ (.A1(_01678_),
    .A2(_05562_),
    .B(_05575_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11544_ (.A1(net23),
    .A2(_05566_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11545_ (.A1(_05561_),
    .A2(_05576_),
    .B(_05577_),
    .C(_05568_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11546_ (.I(\as2650.r123[3][0] ),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11547_ (.I(_05578_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11548_ (.I(\as2650.r123[3][1] ),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11549_ (.I(_05579_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11550_ (.I(\as2650.r123[3][2] ),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11551_ (.I(_05580_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11552_ (.I(\as2650.r123[3][3] ),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11553_ (.I(_05581_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11554_ (.I(\as2650.r123[3][4] ),
    .Z(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11555_ (.I(_05582_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11556_ (.I(\as2650.r123[3][5] ),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11557_ (.I(_05583_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11558_ (.I(\as2650.r123[3][6] ),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11559_ (.I(_05584_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11560_ (.I(\as2650.r123[3][7] ),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11561_ (.I(_05585_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11562_ (.A1(_04517_),
    .A2(_00775_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11563_ (.A1(_00571_),
    .A2(_04535_),
    .B(_05586_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11564_ (.A1(_05292_),
    .A2(_00775_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11565_ (.A1(_00826_),
    .A2(_04535_),
    .B(_05587_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11566_ (.A1(_01711_),
    .A2(_02836_),
    .B(_01280_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11567_ (.A1(_01701_),
    .A2(_01708_),
    .B(_01703_),
    .C(_01034_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11568_ (.A1(_05588_),
    .A2(_05589_),
    .B(_00736_),
    .C(_01078_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11569_ (.A1(_00941_),
    .A2(_05131_),
    .B1(_01113_),
    .B2(_04503_),
    .ZN(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11570_ (.A1(_02787_),
    .A2(_02803_),
    .A3(_02809_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11571_ (.A1(_01460_),
    .A2(_02801_),
    .A3(_02777_),
    .ZN(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11572_ (.A1(_02801_),
    .A2(_03758_),
    .A3(_02777_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11573_ (.A1(_02559_),
    .A2(_05593_),
    .A3(_02796_),
    .A4(_05594_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11574_ (.I(_05189_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11575_ (.A1(_00949_),
    .A2(_05596_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11576_ (.A1(_02781_),
    .A2(_02816_),
    .A3(_05595_),
    .A4(_05597_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11577_ (.A1(_01055_),
    .A2(_03702_),
    .B(_00735_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11578_ (.A1(_00902_),
    .A2(_04567_),
    .B(_05599_),
    .C(_02860_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11579_ (.A1(_02519_),
    .A2(_01529_),
    .A3(_02817_),
    .A4(_05191_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11580_ (.A1(_05598_),
    .A2(_05600_),
    .A3(_05601_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11581_ (.A1(_01107_),
    .A2(_05591_),
    .B(_05592_),
    .C(_05602_),
    .ZN(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11582_ (.A1(_02857_),
    .A2(_04941_),
    .B(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11583_ (.I(_04582_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11584_ (.I(_02546_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11585_ (.A1(_05606_),
    .A2(_04499_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11586_ (.A1(_00626_),
    .A2(_04500_),
    .A3(_05607_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11587_ (.A1(_01217_),
    .A2(_05284_),
    .B1(_02957_),
    .B2(_05388_),
    .C(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11588_ (.A1(_00799_),
    .A2(_05605_),
    .B1(_05609_),
    .B2(_02858_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11589_ (.A1(_05590_),
    .A2(_05604_),
    .A3(_05610_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11590_ (.A1(net78),
    .A2(_05604_),
    .B(_05408_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11591_ (.A1(_05611_),
    .A2(_05612_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11592_ (.I(_02802_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11593_ (.A1(_05292_),
    .A2(_00690_),
    .A3(_05613_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11594_ (.A1(_05460_),
    .A2(_05614_),
    .Z(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11595_ (.A1(_00760_),
    .A2(_01011_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11596_ (.A1(_01778_),
    .A2(_02071_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11597_ (.A1(_01780_),
    .A2(_05617_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11598_ (.A1(_01762_),
    .A2(_05137_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11599_ (.A1(_05146_),
    .A2(_05619_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11600_ (.A1(_02586_),
    .A2(_02585_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11601_ (.A1(_02821_),
    .A2(_02573_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11602_ (.A1(_02132_),
    .A2(_00924_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11603_ (.A1(_00924_),
    .A2(_05618_),
    .B(_05623_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11604_ (.A1(_02872_),
    .A2(_05621_),
    .B1(_05622_),
    .B2(_05624_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11605_ (.A1(_02852_),
    .A2(_02574_),
    .B(_00879_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11606_ (.A1(_00879_),
    .A2(_05625_),
    .B1(_05626_),
    .B2(_01953_),
    .C(_00942_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11607_ (.A1(_05357_),
    .A2(_05620_),
    .B(_05627_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11608_ (.A1(_05616_),
    .A2(_05618_),
    .B1(_05628_),
    .B2(_03840_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11609_ (.A1(_05615_),
    .A2(_05629_),
    .ZN(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11610_ (.A1(_02477_),
    .A2(_05615_),
    .B(_05630_),
    .C(_00745_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11611_ (.A1(_02868_),
    .A2(_00690_),
    .A3(_02802_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11612_ (.A1(_05459_),
    .A2(_05631_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11613_ (.A1(_02703_),
    .A2(_02323_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11614_ (.A1(_05617_),
    .A2(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11615_ (.A1(_01762_),
    .A2(_05138_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11616_ (.A1(_01246_),
    .A2(_00923_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11617_ (.A1(_00924_),
    .A2(_05634_),
    .B(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11618_ (.A1(_02867_),
    .A2(_05621_),
    .B1(_05622_),
    .B2(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11619_ (.A1(_02082_),
    .A2(_05626_),
    .B1(_05638_),
    .B2(_00879_),
    .C(_00942_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11620_ (.A1(_05357_),
    .A2(_05635_),
    .B(_05639_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11621_ (.A1(_05616_),
    .A2(_05634_),
    .B1(_05640_),
    .B2(_04014_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11622_ (.A1(_05632_),
    .A2(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11623_ (.A1(_02703_),
    .A2(_05632_),
    .B(_05642_),
    .C(_00745_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11624_ (.A1(_04537_),
    .A2(_00690_),
    .A3(_05613_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11625_ (.A1(_05460_),
    .A2(_05643_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11626_ (.A1(_01770_),
    .A2(_02324_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11627_ (.A1(_02865_),
    .A2(_05441_),
    .B(_04503_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11628_ (.A1(_01850_),
    .A2(_05645_),
    .B(_05622_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11629_ (.A1(_01240_),
    .A2(_01850_),
    .B(_05647_),
    .ZN(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11630_ (.A1(_05646_),
    .A2(_05648_),
    .B(_04565_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11631_ (.A1(_05645_),
    .A2(_05626_),
    .B(_05649_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11632_ (.A1(_02202_),
    .A2(_05314_),
    .B1(_00942_),
    .B2(_05650_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11633_ (.A1(_05645_),
    .A2(_05616_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11634_ (.A1(_04195_),
    .A2(_05651_),
    .B(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11635_ (.A1(_02202_),
    .A2(_05644_),
    .B(_04381_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11636_ (.A1(_05644_),
    .A2(_05653_),
    .B(_05654_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11637_ (.A1(_01280_),
    .A2(_01446_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11638_ (.A1(_01455_),
    .A2(_05655_),
    .B(_00678_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11639_ (.A1(_01456_),
    .A2(_05655_),
    .B(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11640_ (.A1(_02857_),
    .A2(_02592_),
    .B(_05603_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11641_ (.A1(_02546_),
    .A2(_04521_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11642_ (.A1(_00626_),
    .A2(_04522_),
    .A3(_05659_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11643_ (.A1(_02886_),
    .A2(_05284_),
    .B1(_02957_),
    .B2(_01497_),
    .C(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11644_ (.A1(_00799_),
    .A2(_04857_),
    .B1(_05661_),
    .B2(_02858_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11645_ (.A1(_05657_),
    .A2(_05658_),
    .A3(_05662_),
    .Z(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11646_ (.A1(net52),
    .A2(_05658_),
    .B(_05408_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11647_ (.A1(_05663_),
    .A2(_05664_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11648_ (.A1(_01703_),
    .A2(_02928_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11649_ (.A1(_01701_),
    .A2(_02928_),
    .B(_05665_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11650_ (.A1(_01012_),
    .A2(_02810_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11651_ (.A1(_02856_),
    .A2(_04510_),
    .B(_05667_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11652_ (.A1(_05602_),
    .A2(_05668_),
    .Z(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11653_ (.A1(_02588_),
    .A2(_02962_),
    .B(_04511_),
    .C(_02857_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11654_ (.A1(_05202_),
    .A2(_04720_),
    .B(_05669_),
    .C(_05670_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11655_ (.A1(_00736_),
    .A2(_05666_),
    .B(_05671_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11656_ (.A1(net49),
    .A2(_05669_),
    .B(_05408_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11657_ (.A1(_05672_),
    .A2(_05673_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11658_ (.A1(_02860_),
    .A2(_00677_),
    .A3(_00632_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11659_ (.A1(_05598_),
    .A2(_05601_),
    .A3(_05667_),
    .A4(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11660_ (.A1(_00799_),
    .A2(_00541_),
    .A3(_04517_),
    .B(_05675_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11661_ (.A1(_03233_),
    .A2(_05676_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11662_ (.A1(_05606_),
    .A2(_04518_),
    .B(_04516_),
    .C(_05202_),
    .ZN(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11663_ (.A1(_02933_),
    .A2(_04809_),
    .ZN(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11664_ (.A1(_05675_),
    .A2(_05678_),
    .A3(_05679_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11665_ (.A1(_05677_),
    .A2(_05680_),
    .B(_00755_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11666_ (.A1(_05292_),
    .A2(_05613_),
    .B(_05675_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11667_ (.A1(_05606_),
    .A2(_04513_),
    .B(_04480_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11668_ (.A1(_05314_),
    .A2(_04741_),
    .B1(_05682_),
    .B2(_04514_),
    .C(_05681_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11669_ (.A1(_01862_),
    .A2(_05681_),
    .B(_05683_),
    .C(_00745_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11670_ (.A1(_05606_),
    .A2(_04504_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11671_ (.A1(_05357_),
    .A2(_04505_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11672_ (.A1(_05241_),
    .A2(_04661_),
    .B1(_05684_),
    .B2(_05685_),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11673_ (.A1(_04537_),
    .A2(_05613_),
    .B(_05675_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11674_ (.I0(_05686_),
    .I1(net79),
    .S(_05687_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11675_ (.A1(_00830_),
    .A2(_05688_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11676_ (.I(_05689_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11677_ (.A1(_02854_),
    .A2(_04524_),
    .B(_02362_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11678_ (.A1(_02585_),
    .A2(_04525_),
    .B(_04526_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11679_ (.A1(_05690_),
    .A2(_05691_),
    .B(_00829_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11680_ (.A1(_02977_),
    .A2(_05690_),
    .B(_05692_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11681_ (.A1(_02854_),
    .A2(_04517_),
    .B(_02362_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11682_ (.A1(_02585_),
    .A2(_04518_),
    .B(_04516_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11683_ (.A1(_05693_),
    .A2(_05694_),
    .B(_00829_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11684_ (.A1(_05321_),
    .A2(_05693_),
    .B(_05695_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00014_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00015_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00016_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00017_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00018_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00019_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00020_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00021_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00022_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00023_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00024_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00025_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11697_ (.D(_00026_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00027_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00028_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00029_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00030_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00031_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00032_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00033_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00034_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00035_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00036_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00037_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00038_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00039_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00040_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00041_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00042_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00043_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00044_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00045_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00046_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00047_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00048_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00049_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00050_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00051_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00052_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11724_ (.D(_00053_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00054_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00055_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00056_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00057_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00058_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00059_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11731_ (.D(_00060_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11732_ (.D(_00061_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11733_ (.D(_00062_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00063_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00064_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00065_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00066_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00067_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00068_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00069_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00070_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00071_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00072_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00073_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11745_ (.D(_00074_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00075_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11747_ (.D(_00076_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00077_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00078_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00079_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00080_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00081_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00082_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00083_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00084_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00085_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00086_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00087_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00088_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00089_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11761_ (.D(_00090_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11762_ (.D(_00091_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11763_ (.D(_00092_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11764_ (.D(_00093_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11765_ (.D(_00094_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00095_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11767_ (.D(_00096_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11768_ (.D(_00097_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00098_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00099_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00100_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00101_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00102_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00103_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00104_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00105_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00106_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00107_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00108_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00109_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00110_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00111_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00112_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00113_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00114_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00115_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00116_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00117_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00118_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11790_ (.D(_00119_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00120_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00121_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00122_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00123_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00124_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00125_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00126_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11798_ (.D(_00127_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00128_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00129_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00130_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00131_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00132_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00133_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11805_ (.D(_00134_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11806_ (.D(_00135_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11807_ (.D(_00136_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00137_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00138_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00139_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00140_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11812_ (.D(_00141_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11813_ (.D(_00142_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00143_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00144_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11816_ (.D(_00145_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11817_ (.D(_00146_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11818_ (.D(_00147_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00148_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11820_ (.D(_00149_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11821_ (.D(_00150_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00151_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00152_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00153_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00154_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00155_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00156_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00157_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00158_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00159_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00160_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00161_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00162_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00163_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00164_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00165_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00166_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00167_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00168_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00169_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00170_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00171_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00172_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00173_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00174_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00175_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00176_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11848_ (.D(_00177_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11849_ (.D(_00178_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00179_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00180_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00181_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00182_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00183_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00184_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00185_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00186_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00187_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11859_ (.D(_00188_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00189_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00190_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11862_ (.D(_00191_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00192_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00193_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00194_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00195_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00196_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00197_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00198_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00199_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00200_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00201_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00202_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00203_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00204_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00205_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00206_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00207_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00208_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00209_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00210_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00211_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00212_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00213_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00214_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00215_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00216_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00217_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00218_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00219_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00220_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00221_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00222_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00223_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00224_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00225_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00226_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00227_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00228_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00229_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00230_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00231_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00232_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00233_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00234_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00000_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00005_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00006_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00007_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00008_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00009_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11912_ (.D(_00010_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00011_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00012_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11915_ (.D(_00013_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00001_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00002_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00003_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.cycle[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11919_ (.D(_00004_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00235_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00236_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00237_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00238_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00239_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00240_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00241_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00242_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00243_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11929_ (.D(_00244_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00245_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00246_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00247_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00248_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00249_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00250_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11936_ (.D(_00251_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11937_ (.D(_00252_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00253_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00254_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11940_ (.D(_00255_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00256_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11942_ (.D(_00257_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00258_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11944_ (.D(_00259_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11945_ (.D(_00260_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00261_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00262_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11948_ (.D(_00263_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00264_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11950_ (.D(_00265_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11951_ (.D(_00266_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00267_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00268_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00269_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00270_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00271_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00272_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00273_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00274_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00275_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00276_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00277_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00278_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00279_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.ivec[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00280_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00281_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00282_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00283_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11969_ (.D(_00284_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00285_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00286_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11972_ (.D(_00287_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11973_ (.D(_00288_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11974_ (.D(_00289_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00290_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11976_ (.D(_00291_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11977_ (.D(_00292_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11978_ (.D(_00293_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11979_ (.D(_00294_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11980_ (.D(_00295_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11981_ (.D(_00296_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11982_ (.D(_00297_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11983_ (.D(_00298_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11984_ (.D(_00299_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11985_ (.D(_00300_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11986_ (.D(_00301_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11987_ (.D(_00302_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11988_ (.D(_00303_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11989_ (.D(_00304_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11990_ (.D(_00305_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11991_ (.D(_00306_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11992_ (.D(_00307_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11993_ (.D(_00308_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00309_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00310_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00311_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00312_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00313_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11999_ (.D(_00314_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00315_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00316_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00317_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00318_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12004_ (.D(_00319_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_00320_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00321_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00322_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12008_ (.D(_00323_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00324_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12010_ (.D(_00325_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00326_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00327_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00328_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12014_ (.D(_00329_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12015_ (.D(_00330_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12016_ (.D(_00331_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00332_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00333_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00334_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12020_ (.D(_00335_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12021_ (.D(_00336_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12022_ (.D(_00337_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12023_ (.D(_00338_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12024_ (.D(_00339_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12025_ (.D(_00340_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12026_ (.D(_00341_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12027_ (.D(_00342_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12028_ (.D(_00343_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00344_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12030_ (.D(_00345_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12031_ (.D(_00346_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12032_ (.D(_00347_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12033_ (.D(_00348_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12034_ (.D(_00349_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12035_ (.D(_00350_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00351_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00352_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_00353_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_00354_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_00355_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_00356_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00357_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00358_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00359_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00360_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00361_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00362_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00363_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00364_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00365_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00366_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00367_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(_00368_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(_00369_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(_00370_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(_00371_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(_00372_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(_00373_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(_00374_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(_00375_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_00376_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(_00377_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12063_ (.D(_00378_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_00379_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12065_ (.D(_00380_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12066_ (.D(_00381_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_00382_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00383_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(_00384_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_00385_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(_00386_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_00387_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(_00388_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_00389_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_00390_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00391_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00392_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12078_ (.D(_00393_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(_00394_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(_00395_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(_00396_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(_00397_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(_00398_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(_00399_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(_00400_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(_00401_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(_00402_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(_00403_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(_00404_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(_00405_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12091_ (.D(_00406_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_00407_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00408_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_00409_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_00410_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12096_ (.D(_00411_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12097_ (.D(_00412_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12098_ (.D(_00413_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12099_ (.D(_00414_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12100_ (.D(_00415_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12101_ (.D(_00416_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_00417_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12103_ (.D(_00418_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12104_ (.D(_00419_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12178_ (.I(net82),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12179_ (.I(net82),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12180_ (.I(net82),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12181_ (.I(net82),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12182_ (.I(net83),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12183_ (.I(net83),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12184_ (.I(net83),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12185_ (.I(net29),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout82 (.I(net84),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 fanout85 (.I(net15),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout86 (.I(net79),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout87 (.I(net73),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout88 (.I(net78),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout89 (.I(net48),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout90 (.I(net71),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout91 (.I(net64),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout92 (.I(net56),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout93 (.I(net55),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout94 (.I(net27),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout95 (.I(net28),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout96 (.I(net42),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout97 (.I(net40),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout98 (.I(net33),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout99 (.I(net30),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input10 (.I(io_in[7]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(io_in[8]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input12 (.I(io_in[9]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input6 (.I(io_in[34]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(io_in[35]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input8 (.I(io_in[5]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(io_in[6]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net85),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net30),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net31),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net33),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net34),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output36 (.I(net36),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output37 (.I(net37),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output38 (.I(net38),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output39 (.I(net39),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output40 (.I(net40),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output41 (.I(net41),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output42 (.I(net42),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output43 (.I(net43),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output44 (.I(net44),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output45 (.I(net45),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output46 (.I(net46),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output47 (.I(net47),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output48 (.I(net89),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net53),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net93),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net92),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output57 (.I(net57),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output58 (.I(net58),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output60 (.I(net60),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output61 (.I(net61),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output63 (.I(net63),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net91),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net65),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net67),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net87),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net88),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net86),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire80 (.I(_01079_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire81 (.I(_01268_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_146 (.Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_147 (.Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_148 (.Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_149 (.Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_150 (.Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_151 (.Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_152 (.Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_153 (.Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_154 (.Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_155 (.Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_156 (.Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_157 (.Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_158 (.Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_159 (.Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_160 (.Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_161 (.Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_162 (.Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_163 (.Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_164 (.Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_165 (.Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_166 (.Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_167 (.Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_168 (.Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_169 (.Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_170 (.Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_171 (.Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_172 (.Z(net172));
 assign io_oeb[0] = net146;
 assign io_oeb[13] = net151;
 assign io_oeb[14] = net100;
 assign io_oeb[15] = net101;
 assign io_oeb[16] = net102;
 assign io_oeb[17] = net103;
 assign io_oeb[18] = net104;
 assign io_oeb[19] = net105;
 assign io_oeb[1] = net147;
 assign io_oeb[20] = net106;
 assign io_oeb[21] = net107;
 assign io_oeb[22] = net108;
 assign io_oeb[23] = net109;
 assign io_oeb[24] = net110;
 assign io_oeb[25] = net111;
 assign io_oeb[26] = net112;
 assign io_oeb[27] = net113;
 assign io_oeb[28] = net114;
 assign io_oeb[29] = net115;
 assign io_oeb[2] = net148;
 assign io_oeb[30] = net116;
 assign io_oeb[31] = net117;
 assign io_oeb[32] = net118;
 assign io_oeb[33] = net152;
 assign io_oeb[34] = net153;
 assign io_oeb[35] = net154;
 assign io_oeb[36] = net155;
 assign io_oeb[37] = net156;
 assign io_oeb[3] = net149;
 assign io_oeb[4] = net150;
 assign io_out[0] = net119;
 assign io_out[13] = net124;
 assign io_out[1] = net120;
 assign io_out[2] = net121;
 assign io_out[33] = net125;
 assign io_out[34] = net126;
 assign io_out[35] = net127;
 assign io_out[36] = net128;
 assign io_out[37] = net129;
 assign io_out[3] = net122;
 assign io_out[4] = net123;
 assign la_data_out[32] = net157;
 assign la_data_out[33] = net130;
 assign la_data_out[34] = net158;
 assign la_data_out[35] = net131;
 assign la_data_out[36] = net159;
 assign la_data_out[37] = net132;
 assign la_data_out[38] = net160;
 assign la_data_out[39] = net133;
 assign la_data_out[40] = net161;
 assign la_data_out[41] = net134;
 assign la_data_out[42] = net162;
 assign la_data_out[43] = net135;
 assign la_data_out[44] = net163;
 assign la_data_out[45] = net136;
 assign la_data_out[46] = net164;
 assign la_data_out[47] = net137;
 assign la_data_out[48] = net138;
 assign la_data_out[49] = net165;
 assign la_data_out[50] = net139;
 assign la_data_out[51] = net166;
 assign la_data_out[52] = net140;
 assign la_data_out[53] = net167;
 assign la_data_out[54] = net141;
 assign la_data_out[55] = net168;
 assign la_data_out[56] = net142;
 assign la_data_out[57] = net169;
 assign la_data_out[58] = net143;
 assign la_data_out[59] = net170;
 assign la_data_out[60] = net144;
 assign la_data_out[61] = net171;
 assign la_data_out[62] = net145;
 assign la_data_out[63] = net172;
endmodule

