magic
tech gf180mcuD
magscale 1 10
timestamp 1700712293
<< metal1 >>
rect 1344 51770 53648 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 53648 51770
rect 1344 51684 53648 51718
rect 41246 51602 41298 51614
rect 41246 51538 41298 51550
rect 41470 51602 41522 51614
rect 41470 51538 41522 51550
rect 51214 51378 51266 51390
rect 51214 51314 51266 51326
rect 51438 51378 51490 51390
rect 51438 51314 51490 51326
rect 51662 51378 51714 51390
rect 51662 51314 51714 51326
rect 32398 51266 32450 51278
rect 51326 51266 51378 51278
rect 41906 51214 41918 51266
rect 41970 51214 41982 51266
rect 32398 51202 32450 51214
rect 51326 51202 51378 51214
rect 1344 50986 53648 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 53648 50986
rect 1344 50900 53648 50934
rect 51102 50818 51154 50830
rect 51102 50754 51154 50766
rect 23102 50706 23154 50718
rect 19730 50654 19742 50706
rect 19794 50654 19806 50706
rect 23102 50642 23154 50654
rect 26350 50706 26402 50718
rect 29138 50654 29150 50706
rect 29202 50654 29214 50706
rect 31266 50654 31278 50706
rect 31330 50654 31342 50706
rect 35298 50654 35310 50706
rect 35362 50654 35374 50706
rect 36978 50654 36990 50706
rect 37042 50654 37054 50706
rect 40226 50654 40238 50706
rect 40290 50654 40302 50706
rect 48626 50654 48638 50706
rect 48690 50654 48702 50706
rect 26350 50642 26402 50654
rect 20190 50594 20242 50606
rect 16930 50542 16942 50594
rect 16994 50542 17006 50594
rect 20190 50530 20242 50542
rect 21198 50594 21250 50606
rect 21198 50530 21250 50542
rect 21534 50594 21586 50606
rect 26126 50594 26178 50606
rect 24322 50542 24334 50594
rect 24386 50542 24398 50594
rect 21534 50530 21586 50542
rect 26126 50530 26178 50542
rect 26462 50594 26514 50606
rect 35758 50594 35810 50606
rect 32050 50542 32062 50594
rect 32114 50542 32126 50594
rect 32386 50542 32398 50594
rect 32450 50542 32462 50594
rect 39890 50542 39902 50594
rect 39954 50542 39966 50594
rect 43026 50542 43038 50594
rect 43090 50542 43102 50594
rect 45714 50542 45726 50594
rect 45778 50542 45790 50594
rect 51986 50542 51998 50594
rect 52050 50542 52062 50594
rect 26462 50530 26514 50542
rect 35758 50530 35810 50542
rect 21422 50482 21474 50494
rect 17602 50430 17614 50482
rect 17666 50430 17678 50482
rect 21422 50418 21474 50430
rect 21870 50482 21922 50494
rect 21870 50418 21922 50430
rect 22990 50482 23042 50494
rect 22990 50418 23042 50430
rect 23214 50482 23266 50494
rect 23214 50418 23266 50430
rect 23998 50482 24050 50494
rect 23998 50418 24050 50430
rect 24110 50482 24162 50494
rect 24110 50418 24162 50430
rect 26798 50482 26850 50494
rect 33170 50430 33182 50482
rect 33234 50430 33246 50482
rect 39106 50430 39118 50482
rect 39170 50430 39182 50482
rect 42354 50430 42366 50482
rect 42418 50430 42430 50482
rect 46498 50430 46510 50482
rect 46562 50430 46574 50482
rect 26798 50418 26850 50430
rect 22766 50370 22818 50382
rect 49198 50370 49250 50382
rect 23538 50318 23550 50370
rect 23602 50318 23614 50370
rect 22766 50306 22818 50318
rect 49198 50306 49250 50318
rect 1344 50202 53648 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 53648 50202
rect 1344 50116 53648 50150
rect 20526 50034 20578 50046
rect 20526 49970 20578 49982
rect 21198 50034 21250 50046
rect 21198 49970 21250 49982
rect 21870 50034 21922 50046
rect 21870 49970 21922 49982
rect 26238 50034 26290 50046
rect 26238 49970 26290 49982
rect 33966 50034 34018 50046
rect 33966 49970 34018 49982
rect 36766 50034 36818 50046
rect 36766 49970 36818 49982
rect 37662 50034 37714 50046
rect 37662 49970 37714 49982
rect 41022 50034 41074 50046
rect 41022 49970 41074 49982
rect 49758 50034 49810 50046
rect 49758 49970 49810 49982
rect 49870 50034 49922 50046
rect 49870 49970 49922 49982
rect 49982 50034 50034 50046
rect 49982 49970 50034 49982
rect 21982 49922 22034 49934
rect 21982 49858 22034 49870
rect 23326 49922 23378 49934
rect 23326 49858 23378 49870
rect 23550 49922 23602 49934
rect 23550 49858 23602 49870
rect 25902 49922 25954 49934
rect 25902 49858 25954 49870
rect 26014 49922 26066 49934
rect 26014 49858 26066 49870
rect 27358 49922 27410 49934
rect 27358 49858 27410 49870
rect 27470 49922 27522 49934
rect 27470 49858 27522 49870
rect 33854 49922 33906 49934
rect 33854 49858 33906 49870
rect 37214 49922 37266 49934
rect 37214 49858 37266 49870
rect 37774 49922 37826 49934
rect 37774 49858 37826 49870
rect 41134 49922 41186 49934
rect 48974 49922 49026 49934
rect 43474 49870 43486 49922
rect 43538 49870 43550 49922
rect 51090 49870 51102 49922
rect 51154 49870 51166 49922
rect 41134 49858 41186 49870
rect 48974 49858 49026 49870
rect 19630 49810 19682 49822
rect 19630 49746 19682 49758
rect 19854 49810 19906 49822
rect 19854 49746 19906 49758
rect 21310 49810 21362 49822
rect 21310 49746 21362 49758
rect 26462 49810 26514 49822
rect 26462 49746 26514 49758
rect 26798 49810 26850 49822
rect 26798 49746 26850 49758
rect 26910 49810 26962 49822
rect 26910 49746 26962 49758
rect 27694 49810 27746 49822
rect 33182 49810 33234 49822
rect 34638 49810 34690 49822
rect 32050 49758 32062 49810
rect 32114 49758 32126 49810
rect 34402 49758 34414 49810
rect 34466 49758 34478 49810
rect 27694 49746 27746 49758
rect 33182 49746 33234 49758
rect 34638 49746 34690 49758
rect 34862 49810 34914 49822
rect 36654 49810 36706 49822
rect 35074 49758 35086 49810
rect 35138 49758 35150 49810
rect 34862 49746 34914 49758
rect 36654 49746 36706 49758
rect 36990 49810 37042 49822
rect 39790 49810 39842 49822
rect 39554 49758 39566 49810
rect 39618 49758 39630 49810
rect 36990 49746 37042 49758
rect 39790 49746 39842 49758
rect 40014 49810 40066 49822
rect 42254 49810 42306 49822
rect 48862 49810 48914 49822
rect 40226 49758 40238 49810
rect 40290 49758 40302 49810
rect 42018 49758 42030 49810
rect 42082 49758 42094 49810
rect 42690 49758 42702 49810
rect 42754 49758 42766 49810
rect 49410 49758 49422 49810
rect 49474 49758 49486 49810
rect 50418 49758 50430 49810
rect 50482 49758 50494 49810
rect 40014 49746 40066 49758
rect 42254 49746 42306 49758
rect 48862 49746 48914 49758
rect 26574 49698 26626 49710
rect 23202 49646 23214 49698
rect 23266 49646 23278 49698
rect 26574 49634 26626 49646
rect 28030 49698 28082 49710
rect 36878 49698 36930 49710
rect 29250 49646 29262 49698
rect 29314 49646 29326 49698
rect 31378 49646 31390 49698
rect 31442 49646 31454 49698
rect 34514 49646 34526 49698
rect 34578 49646 34590 49698
rect 28030 49634 28082 49646
rect 36878 49634 36930 49646
rect 37550 49698 37602 49710
rect 37550 49634 37602 49646
rect 39902 49698 39954 49710
rect 39902 49634 39954 49646
rect 40910 49698 40962 49710
rect 45602 49646 45614 49698
rect 45666 49646 45678 49698
rect 53218 49646 53230 49698
rect 53282 49646 53294 49698
rect 40910 49634 40962 49646
rect 20078 49586 20130 49598
rect 20078 49522 20130 49534
rect 21198 49586 21250 49598
rect 21198 49522 21250 49534
rect 21758 49586 21810 49598
rect 21758 49522 21810 49534
rect 34078 49586 34130 49598
rect 34078 49522 34130 49534
rect 42366 49586 42418 49598
rect 42366 49522 42418 49534
rect 48974 49586 49026 49598
rect 48974 49522 49026 49534
rect 1344 49418 53648 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 53648 49418
rect 1344 49332 53648 49366
rect 48750 49250 48802 49262
rect 48750 49186 48802 49198
rect 22094 49138 22146 49150
rect 22094 49074 22146 49086
rect 25678 49138 25730 49150
rect 51886 49138 51938 49150
rect 26450 49086 26462 49138
rect 26514 49086 26526 49138
rect 25678 49074 25730 49086
rect 51886 49074 51938 49086
rect 21646 49026 21698 49038
rect 20738 48974 20750 49026
rect 20802 48974 20814 49026
rect 21646 48962 21698 48974
rect 21758 49026 21810 49038
rect 21758 48962 21810 48974
rect 21982 49026 22034 49038
rect 21982 48962 22034 48974
rect 22654 49026 22706 49038
rect 22654 48962 22706 48974
rect 22990 49026 23042 49038
rect 22990 48962 23042 48974
rect 23438 49026 23490 49038
rect 23438 48962 23490 48974
rect 23662 49026 23714 49038
rect 25566 49026 25618 49038
rect 23986 48974 23998 49026
rect 24050 48974 24062 49026
rect 23662 48962 23714 48974
rect 25566 48962 25618 48974
rect 25790 49026 25842 49038
rect 25790 48962 25842 48974
rect 26014 49026 26066 49038
rect 46062 49026 46114 49038
rect 26338 48974 26350 49026
rect 26402 48974 26414 49026
rect 42690 48974 42702 49026
rect 42754 48974 42766 49026
rect 26014 48962 26066 48974
rect 46062 48962 46114 48974
rect 48974 49026 49026 49038
rect 48974 48962 49026 48974
rect 49198 49026 49250 49038
rect 49634 48974 49646 49026
rect 49698 48974 49710 49026
rect 49198 48962 49250 48974
rect 20414 48914 20466 48926
rect 20414 48850 20466 48862
rect 22430 48914 22482 48926
rect 22430 48850 22482 48862
rect 24558 48914 24610 48926
rect 24558 48850 24610 48862
rect 25342 48914 25394 48926
rect 25342 48850 25394 48862
rect 27134 48914 27186 48926
rect 27134 48850 27186 48862
rect 42254 48914 42306 48926
rect 42254 48850 42306 48862
rect 22766 48802 22818 48814
rect 22766 48738 22818 48750
rect 22878 48802 22930 48814
rect 22878 48738 22930 48750
rect 23550 48802 23602 48814
rect 23550 48738 23602 48750
rect 26574 48802 26626 48814
rect 45950 48802 46002 48814
rect 42466 48750 42478 48802
rect 42530 48750 42542 48802
rect 26574 48738 26626 48750
rect 45950 48738 46002 48750
rect 46398 48802 46450 48814
rect 46398 48738 46450 48750
rect 46622 48802 46674 48814
rect 46622 48738 46674 48750
rect 46734 48802 46786 48814
rect 46734 48738 46786 48750
rect 48302 48802 48354 48814
rect 48302 48738 48354 48750
rect 1344 48634 53648 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 53648 48634
rect 1344 48548 53648 48582
rect 25902 48466 25954 48478
rect 25902 48402 25954 48414
rect 34526 48466 34578 48478
rect 34526 48402 34578 48414
rect 34862 48466 34914 48478
rect 46622 48466 46674 48478
rect 38994 48414 39006 48466
rect 39058 48414 39070 48466
rect 34862 48402 34914 48414
rect 46622 48402 46674 48414
rect 49646 48466 49698 48478
rect 49646 48402 49698 48414
rect 46846 48354 46898 48366
rect 46846 48290 46898 48302
rect 47182 48354 47234 48366
rect 47182 48290 47234 48302
rect 34638 48242 34690 48254
rect 34638 48178 34690 48190
rect 34974 48242 35026 48254
rect 46286 48242 46338 48254
rect 39218 48190 39230 48242
rect 39282 48190 39294 48242
rect 34974 48178 35026 48190
rect 46286 48178 46338 48190
rect 46622 48242 46674 48254
rect 46622 48178 46674 48190
rect 48974 48242 49026 48254
rect 50866 48190 50878 48242
rect 50930 48190 50942 48242
rect 48974 48178 49026 48190
rect 25790 48130 25842 48142
rect 25790 48066 25842 48078
rect 26350 48130 26402 48142
rect 45950 48130 46002 48142
rect 34514 48078 34526 48130
rect 34578 48078 34590 48130
rect 26350 48066 26402 48078
rect 45950 48066 46002 48078
rect 48190 48130 48242 48142
rect 48190 48066 48242 48078
rect 48750 48130 48802 48142
rect 48750 48066 48802 48078
rect 49198 48130 49250 48142
rect 49198 48066 49250 48078
rect 47406 48018 47458 48030
rect 47406 47954 47458 47966
rect 47742 48018 47794 48030
rect 47742 47954 47794 47966
rect 53006 48018 53058 48030
rect 53006 47954 53058 47966
rect 1344 47850 53648 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 53648 47850
rect 1344 47764 53648 47798
rect 27918 47682 27970 47694
rect 27918 47618 27970 47630
rect 37774 47682 37826 47694
rect 37774 47618 37826 47630
rect 12562 47518 12574 47570
rect 12626 47518 12638 47570
rect 19058 47518 19070 47570
rect 19122 47518 19134 47570
rect 34738 47518 34750 47570
rect 34802 47518 34814 47570
rect 42466 47518 42478 47570
rect 42530 47518 42542 47570
rect 49634 47518 49646 47570
rect 49698 47518 49710 47570
rect 51090 47518 51102 47570
rect 51154 47518 51166 47570
rect 20862 47458 20914 47470
rect 9762 47406 9774 47458
rect 9826 47406 9838 47458
rect 16258 47406 16270 47458
rect 16322 47406 16334 47458
rect 20514 47406 20526 47458
rect 20578 47406 20590 47458
rect 20862 47394 20914 47406
rect 21198 47458 21250 47470
rect 21198 47394 21250 47406
rect 21534 47458 21586 47470
rect 42590 47458 42642 47470
rect 28242 47406 28254 47458
rect 28306 47406 28318 47458
rect 31938 47406 31950 47458
rect 32002 47406 32014 47458
rect 39218 47406 39230 47458
rect 39282 47406 39294 47458
rect 42354 47406 42366 47458
rect 42418 47406 42430 47458
rect 21534 47394 21586 47406
rect 42590 47394 42642 47406
rect 42926 47458 42978 47470
rect 42926 47394 42978 47406
rect 49086 47458 49138 47470
rect 49522 47406 49534 47458
rect 49586 47406 49598 47458
rect 49086 47394 49138 47406
rect 20302 47346 20354 47358
rect 10434 47294 10446 47346
rect 10498 47294 10510 47346
rect 16930 47294 16942 47346
rect 16994 47294 17006 47346
rect 20302 47282 20354 47294
rect 21422 47346 21474 47358
rect 21422 47282 21474 47294
rect 21870 47346 21922 47358
rect 21870 47282 21922 47294
rect 24446 47346 24498 47358
rect 24446 47282 24498 47294
rect 24782 47346 24834 47358
rect 35198 47346 35250 47358
rect 37662 47346 37714 47358
rect 25890 47294 25902 47346
rect 25954 47294 25966 47346
rect 32610 47294 32622 47346
rect 32674 47294 32686 47346
rect 36978 47294 36990 47346
rect 37042 47294 37054 47346
rect 24782 47282 24834 47294
rect 35198 47282 35250 47294
rect 37662 47282 37714 47294
rect 37774 47346 37826 47358
rect 37774 47282 37826 47294
rect 38334 47346 38386 47358
rect 48750 47346 48802 47358
rect 39442 47294 39454 47346
rect 39506 47294 39518 47346
rect 38334 47282 38386 47294
rect 48750 47282 48802 47294
rect 50430 47346 50482 47358
rect 50430 47282 50482 47294
rect 50766 47346 50818 47358
rect 50766 47282 50818 47294
rect 9326 47234 9378 47246
rect 9326 47170 9378 47182
rect 19406 47234 19458 47246
rect 20750 47234 20802 47246
rect 19730 47182 19742 47234
rect 19794 47182 19806 47234
rect 19406 47170 19458 47182
rect 20750 47170 20802 47182
rect 26238 47234 26290 47246
rect 26238 47170 26290 47182
rect 28030 47234 28082 47246
rect 31502 47234 31554 47246
rect 31154 47182 31166 47234
rect 31218 47182 31230 47234
rect 28030 47170 28082 47182
rect 31502 47170 31554 47182
rect 37326 47234 37378 47246
rect 37326 47170 37378 47182
rect 42814 47234 42866 47246
rect 42814 47170 42866 47182
rect 46846 47234 46898 47246
rect 46846 47170 46898 47182
rect 48862 47234 48914 47246
rect 48862 47170 48914 47182
rect 50990 47234 51042 47246
rect 50990 47170 51042 47182
rect 1344 47066 53648 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 53648 47066
rect 1344 46980 53648 47014
rect 17950 46898 18002 46910
rect 17950 46834 18002 46846
rect 19294 46898 19346 46910
rect 19294 46834 19346 46846
rect 20974 46898 21026 46910
rect 20974 46834 21026 46846
rect 24110 46898 24162 46910
rect 24110 46834 24162 46846
rect 33182 46898 33234 46910
rect 33182 46834 33234 46846
rect 37102 46898 37154 46910
rect 37102 46834 37154 46846
rect 41806 46898 41858 46910
rect 41806 46834 41858 46846
rect 42142 46898 42194 46910
rect 42142 46834 42194 46846
rect 20526 46786 20578 46798
rect 20526 46722 20578 46734
rect 21086 46786 21138 46798
rect 33406 46786 33458 46798
rect 30034 46734 30046 46786
rect 30098 46734 30110 46786
rect 21086 46722 21138 46734
rect 33406 46722 33458 46734
rect 41582 46786 41634 46798
rect 41582 46722 41634 46734
rect 42926 46786 42978 46798
rect 42926 46722 42978 46734
rect 47854 46786 47906 46798
rect 51090 46734 51102 46786
rect 51154 46734 51166 46786
rect 47854 46722 47906 46734
rect 16158 46674 16210 46686
rect 13010 46622 13022 46674
rect 13074 46622 13086 46674
rect 16158 46610 16210 46622
rect 16382 46674 16434 46686
rect 16382 46610 16434 46622
rect 16606 46674 16658 46686
rect 16606 46610 16658 46622
rect 17502 46674 17554 46686
rect 17502 46610 17554 46622
rect 20638 46674 20690 46686
rect 20638 46610 20690 46622
rect 23102 46674 23154 46686
rect 23102 46610 23154 46622
rect 23214 46674 23266 46686
rect 23214 46610 23266 46622
rect 23326 46674 23378 46686
rect 23326 46610 23378 46622
rect 23774 46674 23826 46686
rect 23774 46610 23826 46622
rect 26238 46674 26290 46686
rect 36430 46674 36482 46686
rect 30706 46622 30718 46674
rect 30770 46622 30782 46674
rect 26238 46610 26290 46622
rect 36430 46610 36482 46622
rect 36878 46674 36930 46686
rect 41246 46674 41298 46686
rect 37426 46622 37438 46674
rect 37490 46622 37502 46674
rect 36878 46610 36930 46622
rect 41246 46610 41298 46622
rect 42030 46674 42082 46686
rect 47742 46674 47794 46686
rect 43362 46622 43374 46674
rect 43426 46622 43438 46674
rect 42030 46610 42082 46622
rect 47742 46610 47794 46622
rect 48078 46674 48130 46686
rect 50418 46622 50430 46674
rect 50482 46622 50494 46674
rect 48078 46610 48130 46622
rect 16270 46562 16322 46574
rect 13682 46510 13694 46562
rect 13746 46510 13758 46562
rect 15810 46510 15822 46562
rect 15874 46510 15886 46562
rect 16270 46498 16322 46510
rect 26798 46562 26850 46574
rect 31278 46562 31330 46574
rect 27906 46510 27918 46562
rect 27970 46510 27982 46562
rect 31154 46510 31166 46562
rect 31218 46510 31230 46562
rect 26798 46498 26850 46510
rect 17390 46450 17442 46462
rect 17390 46386 17442 46398
rect 20526 46450 20578 46462
rect 31169 46447 31215 46510
rect 31278 46498 31330 46510
rect 31726 46562 31778 46574
rect 36206 46562 36258 46574
rect 33058 46510 33070 46562
rect 33122 46510 33134 46562
rect 31726 46498 31778 46510
rect 36206 46498 36258 46510
rect 36990 46562 37042 46574
rect 41918 46562 41970 46574
rect 38210 46510 38222 46562
rect 38274 46510 38286 46562
rect 40338 46510 40350 46562
rect 40402 46510 40414 46562
rect 43026 46510 43038 46562
rect 43090 46510 43102 46562
rect 44146 46510 44158 46562
rect 44210 46510 44222 46562
rect 46274 46510 46286 46562
rect 46338 46510 46350 46562
rect 53218 46510 53230 46562
rect 53282 46510 53294 46562
rect 36990 46498 37042 46510
rect 41918 46498 41970 46510
rect 42702 46450 42754 46462
rect 31826 46447 31838 46450
rect 31169 46401 31838 46447
rect 31826 46398 31838 46401
rect 31890 46398 31902 46450
rect 20526 46386 20578 46398
rect 42702 46386 42754 46398
rect 1344 46282 53648 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 53648 46282
rect 1344 46196 53648 46230
rect 16270 46114 16322 46126
rect 21634 46062 21646 46114
rect 21698 46062 21710 46114
rect 16270 46050 16322 46062
rect 10894 46002 10946 46014
rect 37998 46002 38050 46014
rect 34738 45950 34750 46002
rect 34802 45950 34814 46002
rect 10894 45938 10946 45950
rect 37998 45938 38050 45950
rect 42702 46002 42754 46014
rect 45378 45950 45390 46002
rect 45442 45950 45454 46002
rect 48066 45950 48078 46002
rect 48130 45950 48142 46002
rect 42702 45938 42754 45950
rect 10782 45890 10834 45902
rect 10782 45826 10834 45838
rect 11118 45890 11170 45902
rect 11118 45826 11170 45838
rect 16382 45890 16434 45902
rect 16382 45826 16434 45838
rect 16830 45890 16882 45902
rect 16830 45826 16882 45838
rect 16942 45890 16994 45902
rect 16942 45826 16994 45838
rect 17390 45890 17442 45902
rect 17390 45826 17442 45838
rect 21982 45890 22034 45902
rect 21982 45826 22034 45838
rect 22206 45890 22258 45902
rect 22206 45826 22258 45838
rect 22654 45890 22706 45902
rect 22654 45826 22706 45838
rect 22766 45890 22818 45902
rect 36990 45890 37042 45902
rect 25890 45838 25902 45890
rect 25954 45838 25966 45890
rect 22766 45826 22818 45838
rect 36990 45826 37042 45838
rect 37550 45890 37602 45902
rect 37550 45826 37602 45838
rect 42590 45890 42642 45902
rect 42590 45826 42642 45838
rect 42814 45890 42866 45902
rect 49422 45890 49474 45902
rect 43026 45838 43038 45890
rect 43090 45838 43102 45890
rect 47058 45838 47070 45890
rect 47122 45838 47134 45890
rect 48178 45838 48190 45890
rect 48242 45838 48254 45890
rect 49186 45838 49198 45890
rect 49250 45838 49262 45890
rect 42814 45826 42866 45838
rect 49422 45826 49474 45838
rect 10446 45778 10498 45790
rect 10446 45714 10498 45726
rect 11454 45778 11506 45790
rect 11454 45714 11506 45726
rect 17614 45778 17666 45790
rect 18510 45778 18562 45790
rect 17938 45726 17950 45778
rect 18002 45726 18014 45778
rect 17614 45714 17666 45726
rect 18510 45714 18562 45726
rect 24110 45778 24162 45790
rect 35086 45778 35138 45790
rect 25330 45726 25342 45778
rect 25394 45726 25406 45778
rect 25778 45726 25790 45778
rect 25842 45726 25854 45778
rect 26002 45726 26014 45778
rect 26066 45775 26078 45778
rect 26226 45775 26238 45778
rect 26066 45729 26238 45775
rect 26066 45726 26078 45729
rect 26226 45726 26238 45729
rect 26290 45726 26302 45778
rect 24110 45714 24162 45726
rect 35086 45714 35138 45726
rect 37214 45778 37266 45790
rect 37214 45714 37266 45726
rect 42366 45778 42418 45790
rect 42366 45714 42418 45726
rect 47742 45778 47794 45790
rect 47742 45714 47794 45726
rect 49086 45778 49138 45790
rect 49086 45714 49138 45726
rect 15934 45666 15986 45678
rect 15934 45602 15986 45614
rect 16270 45666 16322 45678
rect 16270 45602 16322 45614
rect 16718 45666 16770 45678
rect 16718 45602 16770 45614
rect 22878 45666 22930 45678
rect 22878 45602 22930 45614
rect 22990 45666 23042 45678
rect 22990 45602 23042 45614
rect 23102 45666 23154 45678
rect 26350 45666 26402 45678
rect 24434 45614 24446 45666
rect 24498 45614 24510 45666
rect 25106 45614 25118 45666
rect 25170 45614 25182 45666
rect 23102 45602 23154 45614
rect 26350 45602 26402 45614
rect 34862 45666 34914 45678
rect 34862 45602 34914 45614
rect 37438 45666 37490 45678
rect 37438 45602 37490 45614
rect 44270 45666 44322 45678
rect 44270 45602 44322 45614
rect 1344 45498 53648 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 53648 45498
rect 1344 45412 53648 45446
rect 11006 45330 11058 45342
rect 11006 45266 11058 45278
rect 14814 45330 14866 45342
rect 14814 45266 14866 45278
rect 17502 45330 17554 45342
rect 17502 45266 17554 45278
rect 23102 45330 23154 45342
rect 23102 45266 23154 45278
rect 23214 45330 23266 45342
rect 23214 45266 23266 45278
rect 24670 45330 24722 45342
rect 24670 45266 24722 45278
rect 41246 45330 41298 45342
rect 41246 45266 41298 45278
rect 41918 45330 41970 45342
rect 41918 45266 41970 45278
rect 48078 45330 48130 45342
rect 48078 45266 48130 45278
rect 48750 45330 48802 45342
rect 48750 45266 48802 45278
rect 12238 45218 12290 45230
rect 42254 45218 42306 45230
rect 12898 45166 12910 45218
rect 12962 45166 12974 45218
rect 19954 45166 19966 45218
rect 20018 45166 20030 45218
rect 28802 45166 28814 45218
rect 28866 45166 28878 45218
rect 33058 45166 33070 45218
rect 33122 45166 33134 45218
rect 38322 45166 38334 45218
rect 38386 45166 38398 45218
rect 38882 45166 38894 45218
rect 38946 45166 38958 45218
rect 12238 45154 12290 45166
rect 42254 45154 42306 45166
rect 42478 45218 42530 45230
rect 42478 45154 42530 45166
rect 43710 45218 43762 45230
rect 43710 45154 43762 45166
rect 48190 45218 48242 45230
rect 48190 45154 48242 45166
rect 48862 45218 48914 45230
rect 48862 45154 48914 45166
rect 10894 45106 10946 45118
rect 10894 45042 10946 45054
rect 11118 45106 11170 45118
rect 11118 45042 11170 45054
rect 11566 45106 11618 45118
rect 11566 45042 11618 45054
rect 11790 45106 11842 45118
rect 11790 45042 11842 45054
rect 12014 45106 12066 45118
rect 12014 45042 12066 45054
rect 12462 45106 12514 45118
rect 14254 45106 14306 45118
rect 13346 45054 13358 45106
rect 13410 45054 13422 45106
rect 13906 45054 13918 45106
rect 13970 45054 13982 45106
rect 12462 45042 12514 45054
rect 14254 45042 14306 45054
rect 17278 45106 17330 45118
rect 17278 45042 17330 45054
rect 17614 45106 17666 45118
rect 21870 45106 21922 45118
rect 29598 45106 29650 45118
rect 32398 45106 32450 45118
rect 41134 45106 41186 45118
rect 18722 45054 18734 45106
rect 18786 45054 18798 45106
rect 19506 45054 19518 45106
rect 19570 45054 19582 45106
rect 20066 45054 20078 45106
rect 20130 45054 20142 45106
rect 22082 45054 22094 45106
rect 22146 45054 22158 45106
rect 25666 45054 25678 45106
rect 25730 45054 25742 45106
rect 29026 45054 29038 45106
rect 29090 45054 29102 45106
rect 31938 45054 31950 45106
rect 32002 45054 32014 45106
rect 33618 45054 33630 45106
rect 33682 45054 33694 45106
rect 34178 45054 34190 45106
rect 34242 45054 34254 45106
rect 37202 45054 37214 45106
rect 37266 45054 37278 45106
rect 38210 45054 38222 45106
rect 38274 45054 38286 45106
rect 46610 45054 46622 45106
rect 46674 45054 46686 45106
rect 47842 45054 47854 45106
rect 47906 45054 47918 45106
rect 50306 45054 50318 45106
rect 50370 45054 50382 45106
rect 17614 45042 17666 45054
rect 21870 45042 21922 45054
rect 29598 45042 29650 45054
rect 32398 45042 32450 45054
rect 41134 45042 41186 45054
rect 14366 44994 14418 45006
rect 22990 44994 23042 45006
rect 31614 44994 31666 45006
rect 34862 44994 34914 45006
rect 39454 44994 39506 45006
rect 12898 44942 12910 44994
rect 12962 44942 12974 44994
rect 22418 44942 22430 44994
rect 22482 44942 22494 44994
rect 26338 44942 26350 44994
rect 26402 44942 26414 44994
rect 28466 44942 28478 44994
rect 28530 44942 28542 44994
rect 33842 44942 33854 44994
rect 33906 44942 33918 44994
rect 35634 44942 35646 44994
rect 35698 44942 35710 44994
rect 14366 44930 14418 44942
rect 22990 44930 23042 44942
rect 31614 44930 31666 44942
rect 34862 44930 34914 44942
rect 39454 44930 39506 44942
rect 42366 44994 42418 45006
rect 47518 44994 47570 45006
rect 45266 44942 45278 44994
rect 45330 44942 45342 44994
rect 42366 44930 42418 44942
rect 47518 44930 47570 44942
rect 49982 44994 50034 45006
rect 51090 44942 51102 44994
rect 51154 44942 51166 44994
rect 53218 44942 53230 44994
rect 53282 44942 53294 44994
rect 49982 44930 50034 44942
rect 12350 44882 12402 44894
rect 41246 44882 41298 44894
rect 19842 44830 19854 44882
rect 19906 44830 19918 44882
rect 22306 44830 22318 44882
rect 22370 44830 22382 44882
rect 12350 44818 12402 44830
rect 41246 44818 41298 44830
rect 1344 44714 53648 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 53648 44714
rect 1344 44628 53648 44662
rect 25902 44546 25954 44558
rect 25902 44482 25954 44494
rect 26238 44546 26290 44558
rect 26238 44482 26290 44494
rect 33294 44546 33346 44558
rect 33294 44482 33346 44494
rect 35534 44546 35586 44558
rect 35534 44482 35586 44494
rect 38446 44546 38498 44558
rect 38446 44482 38498 44494
rect 38894 44546 38946 44558
rect 38894 44482 38946 44494
rect 10110 44434 10162 44446
rect 39454 44434 39506 44446
rect 51774 44434 51826 44446
rect 9650 44382 9662 44434
rect 9714 44382 9726 44434
rect 22082 44382 22094 44434
rect 22146 44382 22158 44434
rect 32050 44382 32062 44434
rect 32114 44382 32126 44434
rect 35074 44382 35086 44434
rect 35138 44382 35150 44434
rect 42130 44382 42142 44434
rect 42194 44382 42206 44434
rect 44258 44382 44270 44434
rect 44322 44382 44334 44434
rect 10110 44370 10162 44382
rect 39454 44370 39506 44382
rect 51774 44370 51826 44382
rect 10670 44322 10722 44334
rect 6850 44270 6862 44322
rect 6914 44270 6926 44322
rect 10670 44258 10722 44270
rect 11342 44322 11394 44334
rect 11342 44258 11394 44270
rect 11790 44322 11842 44334
rect 11790 44258 11842 44270
rect 12574 44322 12626 44334
rect 12574 44258 12626 44270
rect 12686 44322 12738 44334
rect 12686 44258 12738 44270
rect 12798 44322 12850 44334
rect 15934 44322 15986 44334
rect 14466 44270 14478 44322
rect 14530 44270 14542 44322
rect 12798 44258 12850 44270
rect 15934 44258 15986 44270
rect 16494 44322 16546 44334
rect 16494 44258 16546 44270
rect 17278 44322 17330 44334
rect 17278 44258 17330 44270
rect 17502 44322 17554 44334
rect 19742 44322 19794 44334
rect 19282 44270 19294 44322
rect 19346 44270 19358 44322
rect 17502 44258 17554 44270
rect 19742 44258 19794 44270
rect 19966 44322 20018 44334
rect 32398 44322 32450 44334
rect 21298 44270 21310 44322
rect 21362 44270 21374 44322
rect 25106 44270 25118 44322
rect 25170 44270 25182 44322
rect 29250 44270 29262 44322
rect 29314 44270 29326 44322
rect 19966 44258 20018 44270
rect 32398 44258 32450 44270
rect 32622 44322 32674 44334
rect 32622 44258 32674 44270
rect 32846 44322 32898 44334
rect 34078 44322 34130 44334
rect 33618 44270 33630 44322
rect 33682 44270 33694 44322
rect 32846 44258 32898 44270
rect 34078 44258 34130 44270
rect 34750 44322 34802 44334
rect 34750 44258 34802 44270
rect 36094 44322 36146 44334
rect 36094 44258 36146 44270
rect 36318 44322 36370 44334
rect 39006 44322 39058 44334
rect 45054 44322 45106 44334
rect 38546 44270 38558 44322
rect 38610 44270 38622 44322
rect 41346 44270 41358 44322
rect 41410 44270 41422 44322
rect 36318 44258 36370 44270
rect 39006 44258 39058 44270
rect 45054 44258 45106 44270
rect 45614 44322 45666 44334
rect 45614 44258 45666 44270
rect 45950 44322 46002 44334
rect 51102 44322 51154 44334
rect 47506 44270 47518 44322
rect 47570 44270 47582 44322
rect 45950 44258 46002 44270
rect 51102 44258 51154 44270
rect 51214 44322 51266 44334
rect 51214 44258 51266 44270
rect 51662 44322 51714 44334
rect 51662 44258 51714 44270
rect 11678 44210 11730 44222
rect 7522 44158 7534 44210
rect 7586 44158 7598 44210
rect 11678 44146 11730 44158
rect 16046 44210 16098 44222
rect 16046 44146 16098 44158
rect 17838 44210 17890 44222
rect 17838 44146 17890 44158
rect 19854 44210 19906 44222
rect 19854 44146 19906 44158
rect 22542 44210 22594 44222
rect 22542 44146 22594 44158
rect 23998 44210 24050 44222
rect 23998 44146 24050 44158
rect 26126 44210 26178 44222
rect 34414 44210 34466 44222
rect 29922 44158 29934 44210
rect 29986 44158 29998 44210
rect 26126 44146 26178 44158
rect 34414 44146 34466 44158
rect 35758 44210 35810 44222
rect 39790 44210 39842 44222
rect 38210 44158 38222 44210
rect 38274 44158 38286 44210
rect 35758 44146 35810 44158
rect 39790 44146 39842 44158
rect 39902 44210 39954 44222
rect 44942 44210 44994 44222
rect 40674 44158 40686 44210
rect 40738 44158 40750 44210
rect 39902 44146 39954 44158
rect 44942 44146 44994 44158
rect 45502 44210 45554 44222
rect 45502 44146 45554 44158
rect 46062 44210 46114 44222
rect 46062 44146 46114 44158
rect 10782 44098 10834 44110
rect 10782 44034 10834 44046
rect 10894 44098 10946 44110
rect 10894 44034 10946 44046
rect 11454 44098 11506 44110
rect 15150 44098 15202 44110
rect 12114 44046 12126 44098
rect 12178 44046 12190 44098
rect 14690 44046 14702 44098
rect 14754 44046 14766 44098
rect 11454 44034 11506 44046
rect 15150 44034 15202 44046
rect 16158 44098 16210 44110
rect 16158 44034 16210 44046
rect 16830 44098 16882 44110
rect 16830 44034 16882 44046
rect 17390 44098 17442 44110
rect 17390 44034 17442 44046
rect 36430 44098 36482 44110
rect 36430 44034 36482 44046
rect 40126 44098 40178 44110
rect 40126 44034 40178 44046
rect 40350 44098 40402 44110
rect 40350 44034 40402 44046
rect 44718 44098 44770 44110
rect 44718 44034 44770 44046
rect 45278 44098 45330 44110
rect 45278 44034 45330 44046
rect 46286 44098 46338 44110
rect 46286 44034 46338 44046
rect 47742 44098 47794 44110
rect 47742 44034 47794 44046
rect 50878 44098 50930 44110
rect 50878 44034 50930 44046
rect 51326 44098 51378 44110
rect 51326 44034 51378 44046
rect 51886 44098 51938 44110
rect 51886 44034 51938 44046
rect 1344 43930 53648 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 53648 43930
rect 1344 43844 53648 43878
rect 11106 43710 11118 43762
rect 11170 43710 11182 43762
rect 39218 43710 39230 43762
rect 39282 43710 39294 43762
rect 47618 43710 47630 43762
rect 47682 43710 47694 43762
rect 9662 43650 9714 43662
rect 9662 43586 9714 43598
rect 9774 43650 9826 43662
rect 9774 43586 9826 43598
rect 9998 43650 10050 43662
rect 21310 43650 21362 43662
rect 28814 43650 28866 43662
rect 19394 43598 19406 43650
rect 19458 43598 19470 43650
rect 20066 43598 20078 43650
rect 20130 43598 20142 43650
rect 22418 43598 22430 43650
rect 22482 43598 22494 43650
rect 9998 43586 10050 43598
rect 21310 43586 21362 43598
rect 28814 43586 28866 43598
rect 34526 43650 34578 43662
rect 44494 43650 44546 43662
rect 37874 43598 37886 43650
rect 37938 43598 37950 43650
rect 39442 43598 39454 43650
rect 39506 43598 39518 43650
rect 34526 43586 34578 43598
rect 44494 43586 44546 43598
rect 10222 43538 10274 43550
rect 16494 43538 16546 43550
rect 10882 43486 10894 43538
rect 10946 43486 10958 43538
rect 16258 43486 16270 43538
rect 16322 43486 16334 43538
rect 10222 43474 10274 43486
rect 16494 43474 16546 43486
rect 19742 43538 19794 43550
rect 19742 43474 19794 43486
rect 20414 43538 20466 43550
rect 20414 43474 20466 43486
rect 21646 43538 21698 43550
rect 21646 43474 21698 43486
rect 22766 43538 22818 43550
rect 22766 43474 22818 43486
rect 32286 43538 32338 43550
rect 32286 43474 32338 43486
rect 33070 43538 33122 43550
rect 40014 43538 40066 43550
rect 34178 43486 34190 43538
rect 34242 43486 34254 43538
rect 34850 43486 34862 43538
rect 34914 43486 34926 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 38770 43486 38782 43538
rect 38834 43486 38846 43538
rect 33070 43474 33122 43486
rect 40014 43474 40066 43486
rect 41470 43538 41522 43550
rect 41470 43474 41522 43486
rect 47294 43538 47346 43550
rect 51090 43486 51102 43538
rect 51154 43486 51166 43538
rect 47294 43474 47346 43486
rect 17614 43426 17666 43438
rect 17614 43362 17666 43374
rect 31502 43426 31554 43438
rect 31502 43362 31554 43374
rect 32398 43426 32450 43438
rect 39790 43426 39842 43438
rect 33506 43374 33518 43426
rect 33570 43374 33582 43426
rect 35970 43374 35982 43426
rect 36034 43374 36046 43426
rect 32398 43362 32450 43374
rect 39790 43362 39842 43374
rect 41134 43426 41186 43438
rect 46846 43426 46898 43438
rect 41906 43374 41918 43426
rect 41970 43374 41982 43426
rect 41134 43362 41186 43374
rect 46846 43362 46898 43374
rect 47070 43426 47122 43438
rect 47070 43362 47122 43374
rect 53006 43426 53058 43438
rect 53006 43362 53058 43374
rect 16718 43314 16770 43326
rect 16718 43250 16770 43262
rect 16830 43314 16882 43326
rect 16830 43250 16882 43262
rect 31950 43314 32002 43326
rect 31950 43250 32002 43262
rect 32062 43314 32114 43326
rect 32062 43250 32114 43262
rect 34190 43314 34242 43326
rect 40338 43262 40350 43314
rect 40402 43262 40414 43314
rect 34190 43250 34242 43262
rect 1344 43146 53648 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 53648 43146
rect 1344 43060 53648 43094
rect 23550 42978 23602 42990
rect 23550 42914 23602 42926
rect 33742 42978 33794 42990
rect 34066 42926 34078 42978
rect 34130 42975 34142 42978
rect 34850 42975 34862 42978
rect 34130 42929 34862 42975
rect 34130 42926 34142 42929
rect 34850 42926 34862 42929
rect 34914 42926 34926 42978
rect 33742 42914 33794 42926
rect 18062 42866 18114 42878
rect 15474 42814 15486 42866
rect 15538 42814 15550 42866
rect 17602 42814 17614 42866
rect 17666 42814 17678 42866
rect 18062 42802 18114 42814
rect 25454 42866 25506 42878
rect 25454 42802 25506 42814
rect 26350 42866 26402 42878
rect 32398 42866 32450 42878
rect 26674 42814 26686 42866
rect 26738 42814 26750 42866
rect 26350 42802 26402 42814
rect 32398 42802 32450 42814
rect 32734 42866 32786 42878
rect 32734 42802 32786 42814
rect 33854 42866 33906 42878
rect 33854 42802 33906 42814
rect 46734 42866 46786 42878
rect 47842 42814 47854 42866
rect 47906 42814 47918 42866
rect 49970 42814 49982 42866
rect 50034 42814 50046 42866
rect 50978 42814 50990 42866
rect 51042 42814 51054 42866
rect 46734 42802 46786 42814
rect 12462 42754 12514 42766
rect 19182 42754 19234 42766
rect 14802 42702 14814 42754
rect 14866 42702 14878 42754
rect 12462 42690 12514 42702
rect 19182 42690 19234 42702
rect 23662 42754 23714 42766
rect 24110 42754 24162 42766
rect 23874 42702 23886 42754
rect 23938 42702 23950 42754
rect 23662 42690 23714 42702
rect 24110 42690 24162 42702
rect 25006 42754 25058 42766
rect 25006 42690 25058 42702
rect 27918 42754 27970 42766
rect 29262 42754 29314 42766
rect 28354 42702 28366 42754
rect 28418 42702 28430 42754
rect 27918 42690 27970 42702
rect 29262 42690 29314 42702
rect 29486 42754 29538 42766
rect 38558 42754 38610 42766
rect 29698 42702 29710 42754
rect 29762 42702 29774 42754
rect 29486 42690 29538 42702
rect 38558 42690 38610 42702
rect 40014 42754 40066 42766
rect 47058 42702 47070 42754
rect 47122 42702 47134 42754
rect 40014 42690 40066 42702
rect 19070 42642 19122 42654
rect 19070 42578 19122 42590
rect 24446 42642 24498 42654
rect 24446 42578 24498 42590
rect 25230 42642 25282 42654
rect 25230 42578 25282 42590
rect 25566 42642 25618 42654
rect 25566 42578 25618 42590
rect 26014 42642 26066 42654
rect 26014 42578 26066 42590
rect 26574 42642 26626 42654
rect 26574 42578 26626 42590
rect 35870 42642 35922 42654
rect 35870 42578 35922 42590
rect 35982 42642 36034 42654
rect 35982 42578 36034 42590
rect 39902 42642 39954 42654
rect 39902 42578 39954 42590
rect 50654 42642 50706 42654
rect 50654 42578 50706 42590
rect 50878 42642 50930 42654
rect 50878 42578 50930 42590
rect 10446 42530 10498 42542
rect 10446 42466 10498 42478
rect 10894 42530 10946 42542
rect 10894 42466 10946 42478
rect 12574 42530 12626 42542
rect 12574 42466 12626 42478
rect 12798 42530 12850 42542
rect 12798 42466 12850 42478
rect 18846 42530 18898 42542
rect 18846 42466 18898 42478
rect 24670 42530 24722 42542
rect 24670 42466 24722 42478
rect 24782 42530 24834 42542
rect 24782 42466 24834 42478
rect 27470 42530 27522 42542
rect 29598 42530 29650 42542
rect 28578 42478 28590 42530
rect 28642 42478 28654 42530
rect 27470 42466 27522 42478
rect 29598 42466 29650 42478
rect 34414 42530 34466 42542
rect 34414 42466 34466 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 36206 42530 36258 42542
rect 39678 42530 39730 42542
rect 38210 42478 38222 42530
rect 38274 42478 38286 42530
rect 36206 42466 36258 42478
rect 39678 42466 39730 42478
rect 1344 42362 53648 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 53648 42362
rect 1344 42276 53648 42310
rect 11678 42194 11730 42206
rect 13246 42194 13298 42206
rect 24670 42194 24722 42206
rect 12674 42142 12686 42194
rect 12738 42142 12750 42194
rect 23874 42142 23886 42194
rect 23938 42142 23950 42194
rect 11678 42130 11730 42142
rect 13246 42130 13298 42142
rect 24670 42130 24722 42142
rect 25566 42194 25618 42206
rect 25566 42130 25618 42142
rect 25790 42194 25842 42206
rect 25790 42130 25842 42142
rect 34414 42194 34466 42206
rect 34414 42130 34466 42142
rect 34974 42194 35026 42206
rect 34974 42130 35026 42142
rect 49758 42194 49810 42206
rect 49758 42130 49810 42142
rect 10894 42082 10946 42094
rect 10894 42018 10946 42030
rect 11118 42082 11170 42094
rect 11118 42018 11170 42030
rect 11230 42082 11282 42094
rect 11230 42018 11282 42030
rect 13022 42082 13074 42094
rect 33406 42082 33458 42094
rect 27010 42030 27022 42082
rect 27074 42030 27086 42082
rect 13022 42018 13074 42030
rect 33406 42018 33458 42030
rect 33518 42082 33570 42094
rect 33518 42018 33570 42030
rect 34526 42082 34578 42094
rect 34526 42018 34578 42030
rect 35086 42082 35138 42094
rect 35086 42018 35138 42030
rect 41246 42082 41298 42094
rect 41246 42018 41298 42030
rect 49982 42082 50034 42094
rect 51090 42030 51102 42082
rect 51154 42030 51166 42082
rect 49982 42018 50034 42030
rect 10222 41970 10274 41982
rect 10222 41906 10274 41918
rect 10446 41970 10498 41982
rect 10446 41906 10498 41918
rect 10782 41970 10834 41982
rect 10782 41906 10834 41918
rect 12350 41970 12402 41982
rect 12350 41906 12402 41918
rect 12910 41970 12962 41982
rect 21982 41970 22034 41982
rect 13458 41918 13470 41970
rect 13522 41918 13534 41970
rect 12910 41906 12962 41918
rect 21982 41906 22034 41918
rect 23102 41970 23154 41982
rect 23102 41906 23154 41918
rect 23214 41970 23266 41982
rect 23214 41906 23266 41918
rect 23662 41970 23714 41982
rect 23662 41906 23714 41918
rect 24222 41970 24274 41982
rect 24222 41906 24274 41918
rect 24558 41970 24610 41982
rect 24558 41906 24610 41918
rect 25118 41970 25170 41982
rect 29822 41970 29874 41982
rect 26338 41918 26350 41970
rect 26402 41918 26414 41970
rect 25118 41906 25170 41918
rect 29822 41906 29874 41918
rect 33742 41970 33794 41982
rect 33742 41906 33794 41918
rect 34190 41970 34242 41982
rect 34190 41906 34242 41918
rect 41022 41970 41074 41982
rect 41022 41906 41074 41918
rect 41694 41970 41746 41982
rect 47966 41970 48018 41982
rect 47394 41918 47406 41970
rect 47458 41918 47470 41970
rect 41694 41906 41746 41918
rect 47966 41906 48018 41918
rect 49086 41970 49138 41982
rect 49086 41906 49138 41918
rect 49310 41970 49362 41982
rect 49310 41906 49362 41918
rect 49870 41970 49922 41982
rect 50306 41918 50318 41970
rect 50370 41918 50382 41970
rect 49870 41906 49922 41918
rect 10558 41858 10610 41870
rect 10558 41794 10610 41806
rect 12126 41858 12178 41870
rect 12126 41794 12178 41806
rect 23438 41858 23490 41870
rect 23438 41794 23490 41806
rect 25678 41858 25730 41870
rect 25678 41794 25730 41806
rect 29150 41858 29202 41870
rect 29150 41794 29202 41806
rect 41470 41858 41522 41870
rect 44594 41806 44606 41858
rect 44658 41806 44670 41858
rect 46722 41806 46734 41858
rect 46786 41806 46798 41858
rect 53218 41806 53230 41858
rect 53282 41806 53294 41858
rect 41470 41794 41522 41806
rect 34974 41746 35026 41758
rect 34974 41682 35026 41694
rect 1344 41578 53648 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 53648 41578
rect 1344 41492 53648 41526
rect 22430 41410 22482 41422
rect 14018 41358 14030 41410
rect 14082 41358 14094 41410
rect 22430 41346 22482 41358
rect 14814 41298 14866 41310
rect 26126 41298 26178 41310
rect 38558 41298 38610 41310
rect 43486 41298 43538 41310
rect 8082 41246 8094 41298
rect 8146 41246 8158 41298
rect 10210 41246 10222 41298
rect 10274 41246 10286 41298
rect 20514 41246 20526 41298
rect 20578 41246 20590 41298
rect 33170 41246 33182 41298
rect 33234 41246 33246 41298
rect 40898 41246 40910 41298
rect 40962 41246 40974 41298
rect 43026 41246 43038 41298
rect 43090 41246 43102 41298
rect 14814 41234 14866 41246
rect 26126 41234 26178 41246
rect 38558 41234 38610 41246
rect 43486 41234 43538 41246
rect 48526 41298 48578 41310
rect 48526 41234 48578 41246
rect 51886 41298 51938 41310
rect 51886 41234 51938 41246
rect 12350 41186 12402 41198
rect 13470 41186 13522 41198
rect 17726 41186 17778 41198
rect 18734 41186 18786 41198
rect 7298 41134 7310 41186
rect 7362 41134 7374 41186
rect 10882 41134 10894 41186
rect 10946 41134 10958 41186
rect 12674 41134 12686 41186
rect 12738 41134 12750 41186
rect 13682 41134 13694 41186
rect 13746 41134 13758 41186
rect 14018 41134 14030 41186
rect 14082 41134 14094 41186
rect 18274 41134 18286 41186
rect 18338 41134 18350 41186
rect 12350 41122 12402 41134
rect 13470 41122 13522 41134
rect 17726 41122 17778 41134
rect 18734 41122 18786 41134
rect 18958 41186 19010 41198
rect 20414 41186 20466 41198
rect 22654 41186 22706 41198
rect 33742 41186 33794 41198
rect 19954 41134 19966 41186
rect 20018 41134 20030 41186
rect 20626 41134 20638 41186
rect 20690 41134 20702 41186
rect 21746 41134 21758 41186
rect 21810 41134 21822 41186
rect 22866 41134 22878 41186
rect 22930 41134 22942 41186
rect 30370 41134 30382 41186
rect 30434 41134 30446 41186
rect 18958 41122 19010 41134
rect 20414 41122 20466 41134
rect 22654 41122 22706 41134
rect 33742 41122 33794 41134
rect 34078 41186 34130 41198
rect 34078 41122 34130 41134
rect 37102 41186 37154 41198
rect 37102 41122 37154 41134
rect 37214 41186 37266 41198
rect 37214 41122 37266 41134
rect 38110 41186 38162 41198
rect 44382 41186 44434 41198
rect 39666 41134 39678 41186
rect 39730 41134 39742 41186
rect 40114 41134 40126 41186
rect 40178 41134 40190 41186
rect 38110 41122 38162 41134
rect 44382 41122 44434 41134
rect 44718 41186 44770 41198
rect 44718 41122 44770 41134
rect 45166 41186 45218 41198
rect 45166 41122 45218 41134
rect 48862 41186 48914 41198
rect 49970 41134 49982 41186
rect 50034 41134 50046 41186
rect 48862 41122 48914 41134
rect 11118 41074 11170 41086
rect 11118 41010 11170 41022
rect 12910 41074 12962 41086
rect 12910 41010 12962 41022
rect 18062 41074 18114 41086
rect 19182 41074 19234 41086
rect 18498 41022 18510 41074
rect 18562 41022 18574 41074
rect 18062 41010 18114 41022
rect 19182 41010 19234 41022
rect 20190 41074 20242 41086
rect 20190 41010 20242 41022
rect 21198 41074 21250 41086
rect 21198 41010 21250 41022
rect 21310 41074 21362 41086
rect 33854 41074 33906 41086
rect 31042 41022 31054 41074
rect 31106 41022 31118 41074
rect 21310 41010 21362 41022
rect 33854 41010 33906 41022
rect 34302 41074 34354 41086
rect 34302 41010 34354 41022
rect 37550 41074 37602 41086
rect 37550 41010 37602 41022
rect 37774 41074 37826 41086
rect 37774 41010 37826 41022
rect 44046 41074 44098 41086
rect 44046 41010 44098 41022
rect 45390 41074 45442 41086
rect 49186 41022 49198 41074
rect 49250 41022 49262 41074
rect 45390 41010 45442 41022
rect 11566 40962 11618 40974
rect 11566 40898 11618 40910
rect 13022 40962 13074 40974
rect 17838 40962 17890 40974
rect 19630 40962 19682 40974
rect 13906 40910 13918 40962
rect 13970 40910 13982 40962
rect 18610 40910 18622 40962
rect 18674 40910 18686 40962
rect 13022 40898 13074 40910
rect 17838 40898 17890 40910
rect 19630 40898 19682 40910
rect 21534 40962 21586 40974
rect 21534 40898 21586 40910
rect 22766 40962 22818 40974
rect 22766 40898 22818 40910
rect 37326 40962 37378 40974
rect 37326 40898 37378 40910
rect 37998 40962 38050 40974
rect 44158 40962 44210 40974
rect 39442 40910 39454 40962
rect 39506 40910 39518 40962
rect 37998 40898 38050 40910
rect 44158 40898 44210 40910
rect 45054 40962 45106 40974
rect 45054 40898 45106 40910
rect 1344 40794 53648 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 53648 40794
rect 1344 40708 53648 40742
rect 10782 40626 10834 40638
rect 10782 40562 10834 40574
rect 19182 40626 19234 40638
rect 30046 40626 30098 40638
rect 20514 40574 20526 40626
rect 20578 40574 20590 40626
rect 19182 40562 19234 40574
rect 30046 40562 30098 40574
rect 30382 40626 30434 40638
rect 40910 40626 40962 40638
rect 30706 40574 30718 40626
rect 30770 40574 30782 40626
rect 31378 40574 31390 40626
rect 31442 40574 31454 40626
rect 30382 40562 30434 40574
rect 40910 40562 40962 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 33966 40514 34018 40526
rect 21746 40462 21758 40514
rect 21810 40462 21822 40514
rect 22418 40462 22430 40514
rect 22482 40462 22494 40514
rect 33966 40450 34018 40462
rect 34190 40514 34242 40526
rect 41918 40514 41970 40526
rect 36642 40462 36654 40514
rect 36706 40462 36718 40514
rect 41234 40462 41246 40514
rect 41298 40462 41310 40514
rect 34190 40450 34242 40462
rect 41918 40450 41970 40462
rect 19070 40402 19122 40414
rect 23998 40402 24050 40414
rect 20290 40350 20302 40402
rect 20354 40350 20366 40402
rect 20850 40350 20862 40402
rect 20914 40350 20926 40402
rect 19070 40338 19122 40350
rect 23998 40338 24050 40350
rect 31054 40402 31106 40414
rect 31054 40338 31106 40350
rect 33854 40402 33906 40414
rect 33854 40338 33906 40350
rect 34302 40402 34354 40414
rect 42030 40402 42082 40414
rect 35858 40350 35870 40402
rect 35922 40350 35934 40402
rect 34302 40338 34354 40350
rect 42030 40338 42082 40350
rect 44942 40402 44994 40414
rect 44942 40338 44994 40350
rect 45278 40402 45330 40414
rect 45278 40338 45330 40350
rect 45502 40402 45554 40414
rect 50642 40350 50654 40402
rect 50706 40350 50718 40402
rect 45502 40338 45554 40350
rect 14590 40290 14642 40302
rect 33406 40290 33458 40302
rect 39230 40290 39282 40302
rect 21858 40238 21870 40290
rect 21922 40238 21934 40290
rect 38770 40238 38782 40290
rect 38834 40238 38846 40290
rect 14590 40226 14642 40238
rect 33406 40226 33458 40238
rect 39230 40226 39282 40238
rect 45166 40290 45218 40302
rect 45166 40226 45218 40238
rect 53006 40178 53058 40190
rect 14242 40126 14254 40178
rect 14306 40175 14318 40178
rect 14578 40175 14590 40178
rect 14306 40129 14590 40175
rect 14306 40126 14318 40129
rect 14578 40126 14590 40129
rect 14642 40126 14654 40178
rect 53006 40114 53058 40126
rect 1344 40010 53648 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 53648 40010
rect 1344 39924 53648 39958
rect 13918 39842 13970 39854
rect 13918 39778 13970 39790
rect 14590 39842 14642 39854
rect 14590 39778 14642 39790
rect 44942 39842 44994 39854
rect 44942 39778 44994 39790
rect 8990 39730 9042 39742
rect 18958 39730 19010 39742
rect 8530 39678 8542 39730
rect 8594 39678 8606 39730
rect 16146 39678 16158 39730
rect 16210 39678 16222 39730
rect 18386 39678 18398 39730
rect 18450 39678 18462 39730
rect 8990 39666 9042 39678
rect 18958 39666 19010 39678
rect 21646 39730 21698 39742
rect 26350 39730 26402 39742
rect 22754 39678 22766 39730
rect 22818 39678 22830 39730
rect 24882 39678 24894 39730
rect 24946 39678 24958 39730
rect 25890 39678 25902 39730
rect 25954 39727 25966 39730
rect 26114 39727 26126 39730
rect 25954 39681 26126 39727
rect 25954 39678 25966 39681
rect 26114 39678 26126 39681
rect 26178 39678 26190 39730
rect 21646 39666 21698 39678
rect 26350 39666 26402 39678
rect 46062 39730 46114 39742
rect 46386 39678 46398 39730
rect 46450 39678 46462 39730
rect 48514 39678 48526 39730
rect 48578 39678 48590 39730
rect 50866 39678 50878 39730
rect 50930 39678 50942 39730
rect 46062 39666 46114 39678
rect 10558 39618 10610 39630
rect 13806 39618 13858 39630
rect 25230 39618 25282 39630
rect 5730 39566 5742 39618
rect 5794 39566 5806 39618
rect 10098 39566 10110 39618
rect 10162 39566 10174 39618
rect 10994 39566 11006 39618
rect 11058 39566 11070 39618
rect 14242 39566 14254 39618
rect 14306 39566 14318 39618
rect 15474 39566 15486 39618
rect 15538 39566 15550 39618
rect 22082 39566 22094 39618
rect 22146 39566 22158 39618
rect 10558 39554 10610 39566
rect 13806 39554 13858 39566
rect 25230 39554 25282 39566
rect 25566 39618 25618 39630
rect 25566 39554 25618 39566
rect 25790 39618 25842 39630
rect 33518 39618 33570 39630
rect 28130 39566 28142 39618
rect 28194 39566 28206 39618
rect 28354 39566 28366 39618
rect 28418 39566 28430 39618
rect 25790 39554 25842 39566
rect 33518 39554 33570 39566
rect 33854 39618 33906 39630
rect 33854 39554 33906 39566
rect 34190 39618 34242 39630
rect 49186 39566 49198 39618
rect 49250 39566 49262 39618
rect 34190 39554 34242 39566
rect 13470 39506 13522 39518
rect 6402 39454 6414 39506
rect 6466 39454 6478 39506
rect 11218 39454 11230 39506
rect 11282 39454 11294 39506
rect 13470 39442 13522 39454
rect 14702 39506 14754 39518
rect 14702 39442 14754 39454
rect 28590 39506 28642 39518
rect 28590 39442 28642 39454
rect 44830 39506 44882 39518
rect 44830 39442 44882 39454
rect 50542 39506 50594 39518
rect 50542 39442 50594 39454
rect 50766 39506 50818 39518
rect 50766 39442 50818 39454
rect 11678 39394 11730 39406
rect 25342 39394 25394 39406
rect 13906 39342 13918 39394
rect 13970 39342 13982 39394
rect 11678 39330 11730 39342
rect 25342 39330 25394 39342
rect 29262 39394 29314 39406
rect 29262 39330 29314 39342
rect 30718 39394 30770 39406
rect 30718 39330 30770 39342
rect 33630 39394 33682 39406
rect 33630 39330 33682 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 1344 39226 53648 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 53648 39226
rect 1344 39140 53648 39174
rect 6862 39058 6914 39070
rect 6862 38994 6914 39006
rect 10110 39058 10162 39070
rect 10110 38994 10162 39006
rect 10558 39058 10610 39070
rect 10558 38994 10610 39006
rect 15374 39058 15426 39070
rect 15374 38994 15426 39006
rect 17838 39058 17890 39070
rect 17838 38994 17890 39006
rect 24558 39058 24610 39070
rect 24558 38994 24610 39006
rect 29374 39058 29426 39070
rect 29374 38994 29426 39006
rect 33182 39058 33234 39070
rect 33182 38994 33234 39006
rect 41134 39058 41186 39070
rect 41134 38994 41186 39006
rect 44382 39058 44434 39070
rect 44382 38994 44434 39006
rect 49870 39058 49922 39070
rect 49870 38994 49922 39006
rect 49982 39058 50034 39070
rect 49982 38994 50034 39006
rect 29150 38946 29202 38958
rect 40126 38946 40178 38958
rect 9762 38894 9774 38946
rect 9826 38894 9838 38946
rect 12786 38894 12798 38946
rect 12850 38894 12862 38946
rect 18946 38894 18958 38946
rect 19010 38894 19022 38946
rect 30370 38894 30382 38946
rect 30434 38894 30446 38946
rect 29150 38882 29202 38894
rect 40126 38882 40178 38894
rect 40238 38946 40290 38958
rect 40238 38882 40290 38894
rect 41246 38946 41298 38958
rect 41246 38882 41298 38894
rect 44942 38946 44994 38958
rect 44942 38882 44994 38894
rect 45054 38946 45106 38958
rect 51090 38894 51102 38946
rect 51154 38894 51166 38946
rect 45054 38882 45106 38894
rect 6526 38834 6578 38846
rect 6526 38770 6578 38782
rect 6862 38834 6914 38846
rect 6862 38770 6914 38782
rect 7086 38834 7138 38846
rect 23998 38834 24050 38846
rect 12114 38782 12126 38834
rect 12178 38782 12190 38834
rect 18162 38782 18174 38834
rect 18226 38782 18238 38834
rect 7086 38770 7138 38782
rect 23998 38770 24050 38782
rect 27022 38834 27074 38846
rect 29038 38834 29090 38846
rect 40462 38834 40514 38846
rect 27458 38782 27470 38834
rect 27522 38782 27534 38834
rect 29698 38782 29710 38834
rect 29762 38782 29774 38834
rect 35410 38782 35422 38834
rect 35474 38782 35486 38834
rect 27022 38770 27074 38782
rect 29038 38770 29090 38782
rect 40462 38770 40514 38782
rect 40798 38834 40850 38846
rect 40798 38770 40850 38782
rect 41358 38834 41410 38846
rect 41358 38770 41410 38782
rect 44046 38834 44098 38846
rect 44046 38770 44098 38782
rect 44382 38834 44434 38846
rect 44382 38770 44434 38782
rect 44718 38834 44770 38846
rect 44718 38770 44770 38782
rect 49310 38834 49362 38846
rect 49310 38770 49362 38782
rect 49758 38834 49810 38846
rect 50418 38782 50430 38834
rect 50482 38782 50494 38834
rect 49758 38770 49810 38782
rect 27918 38722 27970 38734
rect 14914 38670 14926 38722
rect 14978 38670 14990 38722
rect 21074 38670 21086 38722
rect 21138 38670 21150 38722
rect 27918 38658 27970 38670
rect 28478 38722 28530 38734
rect 38222 38722 38274 38734
rect 32498 38670 32510 38722
rect 32562 38670 32574 38722
rect 36082 38670 36094 38722
rect 36146 38670 36158 38722
rect 28478 38658 28530 38670
rect 38222 38658 38274 38670
rect 38894 38722 38946 38734
rect 53218 38670 53230 38722
rect 53282 38670 53294 38722
rect 38894 38658 38946 38670
rect 45054 38610 45106 38622
rect 45054 38546 45106 38558
rect 1344 38442 53648 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 53648 38442
rect 1344 38356 53648 38390
rect 6862 38274 6914 38286
rect 6862 38210 6914 38222
rect 29150 38274 29202 38286
rect 29150 38210 29202 38222
rect 29710 38274 29762 38286
rect 29710 38210 29762 38222
rect 29822 38274 29874 38286
rect 29822 38210 29874 38222
rect 37102 38162 37154 38174
rect 49982 38162 50034 38174
rect 35970 38110 35982 38162
rect 36034 38110 36046 38162
rect 39218 38110 39230 38162
rect 39282 38110 39294 38162
rect 41346 38110 41358 38162
rect 41410 38110 41422 38162
rect 37102 38098 37154 38110
rect 49982 38098 50034 38110
rect 6974 38050 7026 38062
rect 28590 38050 28642 38062
rect 28130 37998 28142 38050
rect 28194 37998 28206 38050
rect 28354 37998 28366 38050
rect 28418 37998 28430 38050
rect 6974 37986 7026 37998
rect 28590 37986 28642 37998
rect 29262 38050 29314 38062
rect 29262 37986 29314 37998
rect 29486 38050 29538 38062
rect 33058 37998 33070 38050
rect 33122 37998 33134 38050
rect 42130 37998 42142 38050
rect 42194 37998 42206 38050
rect 29486 37986 29538 37998
rect 33730 37886 33742 37938
rect 33794 37886 33806 37938
rect 38098 37886 38110 37938
rect 38162 37886 38174 37938
rect 6862 37826 6914 37838
rect 6862 37762 6914 37774
rect 27246 37826 27298 37838
rect 27246 37762 27298 37774
rect 37774 37826 37826 37838
rect 37774 37762 37826 37774
rect 42590 37826 42642 37838
rect 42590 37762 42642 37774
rect 1344 37658 53648 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 53648 37658
rect 1344 37572 53648 37606
rect 19182 37490 19234 37502
rect 19182 37426 19234 37438
rect 46286 37490 46338 37502
rect 46286 37426 46338 37438
rect 49422 37490 49474 37502
rect 49422 37426 49474 37438
rect 49646 37490 49698 37502
rect 49646 37426 49698 37438
rect 5182 37378 5234 37390
rect 5182 37314 5234 37326
rect 7086 37378 7138 37390
rect 7086 37314 7138 37326
rect 7422 37378 7474 37390
rect 7422 37314 7474 37326
rect 18958 37378 19010 37390
rect 18958 37314 19010 37326
rect 19630 37378 19682 37390
rect 29262 37378 29314 37390
rect 26114 37326 26126 37378
rect 26178 37326 26190 37378
rect 43698 37326 43710 37378
rect 43762 37326 43774 37378
rect 19630 37314 19682 37326
rect 29262 37314 29314 37326
rect 5294 37266 5346 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 5294 37202 5346 37214
rect 5630 37266 5682 37278
rect 5630 37202 5682 37214
rect 5854 37266 5906 37278
rect 5854 37202 5906 37214
rect 6190 37266 6242 37278
rect 15374 37266 15426 37278
rect 18846 37266 18898 37278
rect 29150 37266 29202 37278
rect 48190 37266 48242 37278
rect 6626 37214 6638 37266
rect 6690 37214 6702 37266
rect 6850 37214 6862 37266
rect 6914 37214 6926 37266
rect 9538 37214 9550 37266
rect 9602 37214 9614 37266
rect 13682 37214 13694 37266
rect 13746 37214 13758 37266
rect 14914 37214 14926 37266
rect 14978 37214 14990 37266
rect 16146 37214 16158 37266
rect 16210 37214 16222 37266
rect 17826 37214 17838 37266
rect 17890 37214 17902 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 28802 37214 28814 37266
rect 28866 37214 28878 37266
rect 42914 37214 42926 37266
rect 42978 37214 42990 37266
rect 6190 37202 6242 37214
rect 15374 37202 15426 37214
rect 18846 37202 18898 37214
rect 29150 37202 29202 37214
rect 48190 37202 48242 37214
rect 48974 37266 49026 37278
rect 50642 37214 50654 37266
rect 50706 37214 50718 37266
rect 48974 37202 49026 37214
rect 5742 37154 5794 37166
rect 7534 37154 7586 37166
rect 2482 37102 2494 37154
rect 2546 37102 2558 37154
rect 4610 37102 4622 37154
rect 4674 37102 4686 37154
rect 6962 37102 6974 37154
rect 7026 37102 7038 37154
rect 5742 37090 5794 37102
rect 7534 37090 7586 37102
rect 8990 37154 9042 37166
rect 14142 37154 14194 37166
rect 10322 37102 10334 37154
rect 10386 37102 10398 37154
rect 12450 37102 12462 37154
rect 12514 37102 12526 37154
rect 13794 37102 13806 37154
rect 13858 37102 13870 37154
rect 8990 37090 9042 37102
rect 14142 37090 14194 37102
rect 15486 37154 15538 37166
rect 16830 37154 16882 37166
rect 18510 37154 18562 37166
rect 16370 37102 16382 37154
rect 16434 37102 16446 37154
rect 18162 37102 18174 37154
rect 18226 37102 18238 37154
rect 15486 37090 15538 37102
rect 16830 37090 16882 37102
rect 18510 37090 18562 37102
rect 19854 37154 19906 37166
rect 21422 37154 21474 37166
rect 20738 37102 20750 37154
rect 20802 37102 20814 37154
rect 19854 37090 19906 37102
rect 21422 37090 21474 37102
rect 22990 37154 23042 37166
rect 22990 37090 23042 37102
rect 29822 37154 29874 37166
rect 29822 37090 29874 37102
rect 37438 37154 37490 37166
rect 49534 37154 49586 37166
rect 45826 37102 45838 37154
rect 45890 37102 45902 37154
rect 37438 37090 37490 37102
rect 49534 37090 49586 37102
rect 5182 37042 5234 37054
rect 5182 36978 5234 36990
rect 53006 37042 53058 37054
rect 53006 36978 53058 36990
rect 1344 36874 53648 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 53648 36874
rect 1344 36788 53648 36822
rect 5742 36706 5794 36718
rect 5742 36642 5794 36654
rect 23998 36594 24050 36606
rect 45726 36594 45778 36606
rect 9986 36542 9998 36594
rect 10050 36542 10062 36594
rect 17938 36542 17950 36594
rect 18002 36542 18014 36594
rect 25666 36542 25678 36594
rect 25730 36542 25742 36594
rect 47282 36542 47294 36594
rect 47346 36542 47358 36594
rect 49410 36542 49422 36594
rect 49474 36542 49486 36594
rect 23998 36530 24050 36542
rect 45726 36530 45778 36542
rect 5518 36482 5570 36494
rect 5518 36418 5570 36430
rect 15710 36482 15762 36494
rect 22542 36482 22594 36494
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 18274 36430 18286 36482
rect 18338 36430 18350 36482
rect 22082 36430 22094 36482
rect 22146 36430 22158 36482
rect 15710 36418 15762 36430
rect 22542 36418 22594 36430
rect 23102 36482 23154 36494
rect 39118 36482 39170 36494
rect 40574 36482 40626 36494
rect 23538 36430 23550 36482
rect 23602 36430 23614 36482
rect 24882 36430 24894 36482
rect 24946 36430 24958 36482
rect 25330 36430 25342 36482
rect 25394 36430 25406 36482
rect 39330 36430 39342 36482
rect 39394 36430 39406 36482
rect 23102 36418 23154 36430
rect 39118 36418 39170 36430
rect 40574 36418 40626 36430
rect 43710 36482 43762 36494
rect 43710 36418 43762 36430
rect 44830 36482 44882 36494
rect 44830 36418 44882 36430
rect 45502 36482 45554 36494
rect 45502 36418 45554 36430
rect 46174 36482 46226 36494
rect 50990 36482 51042 36494
rect 46498 36430 46510 36482
rect 46562 36430 46574 36482
rect 46174 36418 46226 36430
rect 50990 36418 51042 36430
rect 51214 36482 51266 36494
rect 51214 36418 51266 36430
rect 9550 36370 9602 36382
rect 9550 36306 9602 36318
rect 10222 36370 10274 36382
rect 22654 36370 22706 36382
rect 40686 36370 40738 36382
rect 16594 36318 16606 36370
rect 16658 36318 16670 36370
rect 18162 36318 18174 36370
rect 18226 36318 18238 36370
rect 24322 36318 24334 36370
rect 24386 36318 24398 36370
rect 26002 36318 26014 36370
rect 26066 36318 26078 36370
rect 10222 36306 10274 36318
rect 22654 36306 22706 36318
rect 40686 36306 40738 36318
rect 42254 36370 42306 36382
rect 42254 36306 42306 36318
rect 42366 36370 42418 36382
rect 42366 36306 42418 36318
rect 43822 36370 43874 36382
rect 43822 36306 43874 36318
rect 44942 36370 44994 36382
rect 44942 36306 44994 36318
rect 45950 36370 46002 36382
rect 45950 36306 46002 36318
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 5854 36258 5906 36270
rect 5854 36194 5906 36206
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 9214 36258 9266 36270
rect 9214 36194 9266 36206
rect 9998 36258 10050 36270
rect 9998 36194 10050 36206
rect 10670 36258 10722 36270
rect 10670 36194 10722 36206
rect 38334 36258 38386 36270
rect 38334 36194 38386 36206
rect 38782 36258 38834 36270
rect 38782 36194 38834 36206
rect 38894 36258 38946 36270
rect 38894 36194 38946 36206
rect 39006 36258 39058 36270
rect 39006 36194 39058 36206
rect 40910 36258 40962 36270
rect 40910 36194 40962 36206
rect 42030 36258 42082 36270
rect 42030 36194 42082 36206
rect 42926 36258 42978 36270
rect 42926 36194 42978 36206
rect 44046 36258 44098 36270
rect 44046 36194 44098 36206
rect 45166 36258 45218 36270
rect 45166 36194 45218 36206
rect 50766 36258 50818 36270
rect 50766 36194 50818 36206
rect 51102 36258 51154 36270
rect 51102 36194 51154 36206
rect 1344 36090 53648 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 53648 36090
rect 1344 36004 53648 36038
rect 5294 35922 5346 35934
rect 6862 35922 6914 35934
rect 5730 35870 5742 35922
rect 5794 35870 5806 35922
rect 5294 35858 5346 35870
rect 6862 35858 6914 35870
rect 6974 35922 7026 35934
rect 6974 35858 7026 35870
rect 9998 35922 10050 35934
rect 9998 35858 10050 35870
rect 16606 35922 16658 35934
rect 16606 35858 16658 35870
rect 32622 35922 32674 35934
rect 32622 35858 32674 35870
rect 43038 35922 43090 35934
rect 43038 35858 43090 35870
rect 44158 35922 44210 35934
rect 46174 35922 46226 35934
rect 44370 35870 44382 35922
rect 44434 35870 44446 35922
rect 44158 35858 44210 35870
rect 46174 35858 46226 35870
rect 49982 35922 50034 35934
rect 49982 35858 50034 35870
rect 5182 35810 5234 35822
rect 5182 35746 5234 35758
rect 5406 35810 5458 35822
rect 5406 35746 5458 35758
rect 6302 35810 6354 35822
rect 6302 35746 6354 35758
rect 7310 35810 7362 35822
rect 7310 35746 7362 35758
rect 9550 35810 9602 35822
rect 9550 35746 9602 35758
rect 22878 35810 22930 35822
rect 22878 35746 22930 35758
rect 26238 35810 26290 35822
rect 34078 35810 34130 35822
rect 44830 35810 44882 35822
rect 30594 35758 30606 35810
rect 30658 35758 30670 35810
rect 32386 35758 32398 35810
rect 32450 35758 32462 35810
rect 40898 35758 40910 35810
rect 40962 35758 40974 35810
rect 26238 35746 26290 35758
rect 34078 35746 34130 35758
rect 44830 35746 44882 35758
rect 6190 35698 6242 35710
rect 7086 35698 7138 35710
rect 12126 35698 12178 35710
rect 16046 35698 16098 35710
rect 19742 35698 19794 35710
rect 6514 35646 6526 35698
rect 6578 35646 6590 35698
rect 9762 35646 9774 35698
rect 9826 35646 9838 35698
rect 11778 35646 11790 35698
rect 11842 35646 11854 35698
rect 12898 35646 12910 35698
rect 12962 35646 12974 35698
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 15586 35646 15598 35698
rect 15650 35646 15662 35698
rect 17826 35646 17838 35698
rect 17890 35646 17902 35698
rect 18274 35646 18286 35698
rect 18338 35646 18350 35698
rect 19282 35646 19294 35698
rect 19346 35646 19358 35698
rect 6190 35634 6242 35646
rect 7086 35634 7138 35646
rect 12126 35634 12178 35646
rect 16046 35634 16098 35646
rect 19742 35634 19794 35646
rect 20414 35698 20466 35710
rect 26798 35698 26850 35710
rect 22194 35646 22206 35698
rect 22258 35646 22270 35698
rect 25778 35646 25790 35698
rect 25842 35646 25854 35698
rect 20414 35634 20466 35646
rect 26798 35634 26850 35646
rect 30158 35698 30210 35710
rect 30158 35634 30210 35646
rect 30942 35698 30994 35710
rect 33182 35698 33234 35710
rect 31602 35646 31614 35698
rect 31666 35646 31678 35698
rect 32162 35646 32174 35698
rect 32226 35646 32238 35698
rect 30942 35634 30994 35646
rect 33182 35634 33234 35646
rect 33966 35698 34018 35710
rect 33966 35634 34018 35646
rect 34302 35698 34354 35710
rect 38894 35698 38946 35710
rect 42702 35698 42754 35710
rect 35410 35646 35422 35698
rect 35474 35646 35486 35698
rect 41122 35646 41134 35698
rect 41186 35646 41198 35698
rect 41682 35646 41694 35698
rect 41746 35646 41758 35698
rect 42130 35646 42142 35698
rect 42194 35646 42206 35698
rect 34302 35634 34354 35646
rect 38894 35634 38946 35646
rect 42702 35634 42754 35646
rect 43710 35698 43762 35710
rect 43710 35634 43762 35646
rect 43934 35698 43986 35710
rect 43934 35634 43986 35646
rect 44382 35698 44434 35710
rect 50306 35646 50318 35698
rect 50370 35646 50382 35698
rect 44382 35634 44434 35646
rect 12238 35586 12290 35598
rect 9986 35534 9998 35586
rect 10050 35534 10062 35586
rect 12238 35522 12290 35534
rect 13582 35586 13634 35598
rect 13582 35522 13634 35534
rect 14030 35586 14082 35598
rect 14030 35522 14082 35534
rect 15150 35586 15202 35598
rect 15150 35522 15202 35534
rect 18510 35586 18562 35598
rect 18510 35522 18562 35534
rect 19854 35586 19906 35598
rect 23438 35586 23490 35598
rect 21970 35534 21982 35586
rect 22034 35534 22046 35586
rect 19854 35522 19906 35534
rect 23438 35522 23490 35534
rect 24222 35586 24274 35598
rect 27134 35586 27186 35598
rect 25330 35534 25342 35586
rect 25394 35534 25406 35586
rect 24222 35522 24274 35534
rect 27134 35522 27186 35534
rect 29038 35586 29090 35598
rect 29038 35522 29090 35534
rect 29486 35586 29538 35598
rect 29486 35522 29538 35534
rect 34638 35586 34690 35598
rect 38222 35586 38274 35598
rect 36082 35534 36094 35586
rect 36146 35534 36158 35586
rect 34638 35522 34690 35534
rect 38222 35522 38274 35534
rect 39790 35586 39842 35598
rect 39790 35522 39842 35534
rect 40350 35586 40402 35598
rect 40350 35522 40402 35534
rect 45278 35586 45330 35598
rect 45278 35522 45330 35534
rect 49198 35586 49250 35598
rect 51090 35534 51102 35586
rect 51154 35534 51166 35586
rect 53218 35534 53230 35586
rect 53282 35534 53294 35586
rect 49198 35522 49250 35534
rect 42478 35474 42530 35486
rect 34402 35422 34414 35474
rect 34466 35471 34478 35474
rect 34850 35471 34862 35474
rect 34466 35425 34862 35471
rect 34466 35422 34478 35425
rect 34850 35422 34862 35425
rect 34914 35422 34926 35474
rect 42478 35410 42530 35422
rect 1344 35306 53648 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 53648 35306
rect 1344 35220 53648 35254
rect 33854 35138 33906 35150
rect 33854 35074 33906 35086
rect 36094 35138 36146 35150
rect 36094 35074 36146 35086
rect 50878 35138 50930 35150
rect 50878 35074 50930 35086
rect 5182 35026 5234 35038
rect 10222 35026 10274 35038
rect 4610 34974 4622 35026
rect 4674 34974 4686 35026
rect 8418 34974 8430 35026
rect 8482 34974 8494 35026
rect 5182 34962 5234 34974
rect 10222 34962 10274 34974
rect 11566 35026 11618 35038
rect 11566 34962 11618 34974
rect 12462 35026 12514 35038
rect 30158 35026 30210 35038
rect 38446 35026 38498 35038
rect 17490 34974 17502 35026
rect 17554 34974 17566 35026
rect 31714 34974 31726 35026
rect 31778 34974 31790 35026
rect 35074 34974 35086 35026
rect 35138 34974 35150 35026
rect 12462 34962 12514 34974
rect 30158 34962 30210 34974
rect 38446 34962 38498 34974
rect 40126 35026 40178 35038
rect 40126 34962 40178 34974
rect 45166 35026 45218 35038
rect 46722 34974 46734 35026
rect 46786 34974 46798 35026
rect 48850 34974 48862 35026
rect 48914 34974 48926 35026
rect 51090 34974 51102 35026
rect 51154 34974 51166 35026
rect 45166 34962 45218 34974
rect 10334 34914 10386 34926
rect 19630 34914 19682 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 7522 34862 7534 34914
rect 7586 34862 7598 34914
rect 9874 34862 9886 34914
rect 9938 34862 9950 34914
rect 15698 34862 15710 34914
rect 15762 34862 15774 34914
rect 19058 34862 19070 34914
rect 19122 34862 19134 34914
rect 10334 34850 10386 34862
rect 19630 34850 19682 34862
rect 31054 34914 31106 34926
rect 33630 34914 33682 34926
rect 31938 34862 31950 34914
rect 32002 34862 32014 34914
rect 32610 34862 32622 34914
rect 32674 34862 32686 34914
rect 32946 34862 32958 34914
rect 33010 34862 33022 34914
rect 31054 34850 31106 34862
rect 33630 34850 33682 34862
rect 38894 34914 38946 34926
rect 38894 34850 38946 34862
rect 39230 34914 39282 34926
rect 41582 34914 41634 34926
rect 39778 34862 39790 34914
rect 39842 34862 39854 34914
rect 39230 34850 39282 34862
rect 41582 34850 41634 34862
rect 45278 34914 45330 34926
rect 49534 34914 49586 34926
rect 45938 34862 45950 34914
rect 46002 34862 46014 34914
rect 45278 34850 45330 34862
rect 49534 34850 49586 34862
rect 49758 34914 49810 34926
rect 49758 34850 49810 34862
rect 25342 34802 25394 34814
rect 2482 34750 2494 34802
rect 2546 34750 2558 34802
rect 18498 34750 18510 34802
rect 18562 34750 18574 34802
rect 20066 34750 20078 34802
rect 20130 34750 20142 34802
rect 25342 34738 25394 34750
rect 25678 34802 25730 34814
rect 34750 34802 34802 34814
rect 31266 34750 31278 34802
rect 31330 34750 31342 34802
rect 33394 34750 33406 34802
rect 33458 34750 33470 34802
rect 25678 34738 25730 34750
rect 34750 34738 34802 34750
rect 35534 34802 35586 34814
rect 35534 34738 35586 34750
rect 39454 34802 39506 34814
rect 39454 34738 39506 34750
rect 40462 34802 40514 34814
rect 40462 34738 40514 34750
rect 42478 34802 42530 34814
rect 42478 34738 42530 34750
rect 42590 34802 42642 34814
rect 42590 34738 42642 34750
rect 45054 34802 45106 34814
rect 45054 34738 45106 34750
rect 45614 34802 45666 34814
rect 45614 34738 45666 34750
rect 49646 34802 49698 34814
rect 49646 34738 49698 34750
rect 10110 34690 10162 34702
rect 10110 34626 10162 34638
rect 10446 34690 10498 34702
rect 10446 34626 10498 34638
rect 11006 34690 11058 34702
rect 11006 34626 11058 34638
rect 18174 34690 18226 34702
rect 26126 34690 26178 34702
rect 19170 34638 19182 34690
rect 19234 34638 19246 34690
rect 18174 34626 18226 34638
rect 26126 34626 26178 34638
rect 29710 34690 29762 34702
rect 29710 34626 29762 34638
rect 30606 34690 30658 34702
rect 30606 34626 30658 34638
rect 33966 34690 34018 34702
rect 33966 34626 34018 34638
rect 34190 34690 34242 34702
rect 34190 34626 34242 34638
rect 34974 34690 35026 34702
rect 34974 34626 35026 34638
rect 35198 34690 35250 34702
rect 35198 34626 35250 34638
rect 35758 34690 35810 34702
rect 35758 34626 35810 34638
rect 35982 34690 36034 34702
rect 35982 34626 36034 34638
rect 39006 34690 39058 34702
rect 39006 34626 39058 34638
rect 39118 34690 39170 34702
rect 39118 34626 39170 34638
rect 40014 34690 40066 34702
rect 40014 34626 40066 34638
rect 40238 34690 40290 34702
rect 40238 34626 40290 34638
rect 41022 34690 41074 34702
rect 41022 34626 41074 34638
rect 42142 34690 42194 34702
rect 42142 34626 42194 34638
rect 42814 34690 42866 34702
rect 42814 34626 42866 34638
rect 43374 34690 43426 34702
rect 43374 34626 43426 34638
rect 44382 34690 44434 34702
rect 44382 34626 44434 34638
rect 49310 34690 49362 34702
rect 49310 34626 49362 34638
rect 50654 34690 50706 34702
rect 50654 34626 50706 34638
rect 51102 34690 51154 34702
rect 51102 34626 51154 34638
rect 1344 34522 53648 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 53648 34522
rect 1344 34436 53648 34470
rect 6526 34354 6578 34366
rect 6526 34290 6578 34302
rect 11342 34354 11394 34366
rect 11342 34290 11394 34302
rect 20526 34354 20578 34366
rect 20526 34290 20578 34302
rect 24670 34354 24722 34366
rect 24670 34290 24722 34302
rect 33406 34354 33458 34366
rect 33406 34290 33458 34302
rect 33630 34354 33682 34366
rect 33630 34290 33682 34302
rect 34302 34354 34354 34366
rect 34302 34290 34354 34302
rect 35422 34354 35474 34366
rect 35422 34290 35474 34302
rect 37886 34354 37938 34366
rect 37886 34290 37938 34302
rect 38446 34354 38498 34366
rect 38446 34290 38498 34302
rect 39566 34354 39618 34366
rect 39566 34290 39618 34302
rect 50094 34354 50146 34366
rect 50094 34290 50146 34302
rect 6750 34242 6802 34254
rect 6750 34178 6802 34190
rect 7198 34242 7250 34254
rect 7198 34178 7250 34190
rect 7422 34242 7474 34254
rect 7422 34178 7474 34190
rect 7534 34242 7586 34254
rect 7534 34178 7586 34190
rect 10110 34242 10162 34254
rect 10110 34178 10162 34190
rect 13582 34242 13634 34254
rect 13582 34178 13634 34190
rect 15598 34242 15650 34254
rect 15598 34178 15650 34190
rect 19294 34242 19346 34254
rect 33294 34242 33346 34254
rect 24322 34190 24334 34242
rect 24386 34190 24398 34242
rect 19294 34178 19346 34190
rect 33294 34178 33346 34190
rect 33966 34242 34018 34254
rect 33966 34178 34018 34190
rect 34078 34242 34130 34254
rect 34078 34178 34130 34190
rect 34862 34242 34914 34254
rect 34862 34178 34914 34190
rect 38670 34242 38722 34254
rect 42914 34190 42926 34242
rect 42978 34190 42990 34242
rect 44370 34190 44382 34242
rect 44434 34190 44446 34242
rect 38670 34178 38722 34190
rect 5294 34130 5346 34142
rect 5294 34066 5346 34078
rect 6190 34130 6242 34142
rect 6190 34066 6242 34078
rect 6414 34130 6466 34142
rect 6414 34066 6466 34078
rect 6974 34130 7026 34142
rect 6974 34066 7026 34078
rect 8990 34130 9042 34142
rect 12574 34130 12626 34142
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 8990 34066 9042 34078
rect 12574 34066 12626 34078
rect 12686 34130 12738 34142
rect 19182 34130 19234 34142
rect 34526 34130 34578 34142
rect 38558 34130 38610 34142
rect 49646 34130 49698 34142
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 15026 34078 15038 34130
rect 15090 34078 15102 34130
rect 18610 34078 18622 34130
rect 18674 34078 18686 34130
rect 20850 34078 20862 34130
rect 20914 34078 20926 34130
rect 27122 34078 27134 34130
rect 27186 34078 27198 34130
rect 38210 34078 38222 34130
rect 38274 34078 38286 34130
rect 38882 34078 38894 34130
rect 38946 34078 38958 34130
rect 43026 34078 43038 34130
rect 43090 34078 43102 34130
rect 43810 34078 43822 34130
rect 43874 34078 43886 34130
rect 44146 34078 44158 34130
rect 44210 34078 44222 34130
rect 12686 34066 12738 34078
rect 19182 34066 19234 34078
rect 34526 34066 34578 34078
rect 38558 34066 38610 34078
rect 49646 34066 49698 34078
rect 50318 34130 50370 34142
rect 50642 34078 50654 34130
rect 50706 34078 50718 34130
rect 50318 34066 50370 34078
rect 9998 34018 10050 34030
rect 23774 34018 23826 34030
rect 29934 34018 29986 34030
rect 10882 33966 10894 34018
rect 10946 33966 10958 34018
rect 15586 33966 15598 34018
rect 15650 33966 15662 34018
rect 21634 33966 21646 34018
rect 21698 33966 21710 34018
rect 27794 33966 27806 34018
rect 27858 33966 27870 34018
rect 9998 33954 10050 33966
rect 23774 33954 23826 33966
rect 29934 33954 29986 33966
rect 30606 34018 30658 34030
rect 30606 33954 30658 33966
rect 35758 34018 35810 34030
rect 35758 33954 35810 33966
rect 42590 34018 42642 34030
rect 42590 33954 42642 33966
rect 48862 34018 48914 34030
rect 48862 33954 48914 33966
rect 50206 34018 50258 34030
rect 50206 33954 50258 33966
rect 5518 33906 5570 33918
rect 5518 33842 5570 33854
rect 5742 33906 5794 33918
rect 5742 33842 5794 33854
rect 8878 33906 8930 33918
rect 8878 33842 8930 33854
rect 9662 33906 9714 33918
rect 9662 33842 9714 33854
rect 9774 33906 9826 33918
rect 9774 33842 9826 33854
rect 53006 33906 53058 33918
rect 53006 33842 53058 33854
rect 1344 33738 53648 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 53648 33738
rect 1344 33652 53648 33686
rect 43486 33570 43538 33582
rect 43486 33506 43538 33518
rect 50878 33570 50930 33582
rect 50878 33506 50930 33518
rect 7982 33458 8034 33470
rect 12910 33458 12962 33470
rect 21982 33458 22034 33470
rect 28254 33458 28306 33470
rect 9986 33406 9998 33458
rect 10050 33406 10062 33458
rect 16370 33406 16382 33458
rect 16434 33406 16446 33458
rect 24882 33406 24894 33458
rect 24946 33406 24958 33458
rect 7982 33394 8034 33406
rect 12910 33394 12962 33406
rect 21982 33394 22034 33406
rect 28254 33394 28306 33406
rect 29486 33458 29538 33470
rect 29486 33394 29538 33406
rect 32846 33458 32898 33470
rect 32846 33394 32898 33406
rect 33854 33458 33906 33470
rect 33854 33394 33906 33406
rect 34414 33458 34466 33470
rect 34414 33394 34466 33406
rect 44830 33458 44882 33470
rect 44830 33394 44882 33406
rect 21758 33346 21810 33358
rect 8306 33294 8318 33346
rect 8370 33294 8382 33346
rect 9874 33294 9886 33346
rect 9938 33294 9950 33346
rect 10210 33294 10222 33346
rect 10274 33294 10286 33346
rect 10994 33294 11006 33346
rect 11058 33294 11070 33346
rect 17378 33294 17390 33346
rect 17442 33294 17454 33346
rect 21758 33282 21810 33294
rect 22094 33346 22146 33358
rect 22094 33282 22146 33294
rect 22430 33346 22482 33358
rect 41694 33346 41746 33358
rect 45390 33346 45442 33358
rect 27794 33294 27806 33346
rect 27858 33294 27870 33346
rect 31602 33294 31614 33346
rect 31666 33294 31678 33346
rect 32386 33294 32398 33346
rect 32450 33294 32462 33346
rect 42130 33294 42142 33346
rect 42194 33294 42206 33346
rect 42690 33294 42702 33346
rect 42754 33294 42766 33346
rect 43138 33294 43150 33346
rect 43202 33294 43214 33346
rect 22430 33282 22482 33294
rect 41694 33282 41746 33294
rect 45390 33282 45442 33294
rect 46062 33346 46114 33358
rect 46062 33282 46114 33294
rect 48750 33346 48802 33358
rect 48750 33282 48802 33294
rect 49422 33346 49474 33358
rect 49422 33282 49474 33294
rect 27010 33182 27022 33234
rect 27074 33182 27086 33234
rect 42018 33182 42030 33234
rect 42082 33182 42094 33234
rect 49074 33182 49086 33234
rect 49138 33182 49150 33234
rect 49746 33182 49758 33234
rect 49810 33182 49822 33234
rect 8094 33122 8146 33134
rect 8094 33058 8146 33070
rect 9214 33122 9266 33134
rect 17950 33122 18002 33134
rect 11218 33070 11230 33122
rect 11282 33070 11294 33122
rect 9214 33058 9266 33070
rect 17950 33058 18002 33070
rect 37214 33122 37266 33134
rect 37214 33058 37266 33070
rect 39902 33122 39954 33134
rect 50206 33122 50258 33134
rect 45714 33070 45726 33122
rect 45778 33070 45790 33122
rect 39902 33058 39954 33070
rect 50206 33058 50258 33070
rect 50990 33122 51042 33134
rect 50990 33058 51042 33070
rect 51102 33122 51154 33134
rect 51102 33058 51154 33070
rect 51662 33122 51714 33134
rect 51662 33058 51714 33070
rect 1344 32954 53648 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 53648 32954
rect 1344 32868 53648 32902
rect 9662 32786 9714 32798
rect 9662 32722 9714 32734
rect 21646 32786 21698 32798
rect 21646 32722 21698 32734
rect 25566 32786 25618 32798
rect 25566 32722 25618 32734
rect 26238 32786 26290 32798
rect 26238 32722 26290 32734
rect 33518 32786 33570 32798
rect 37550 32786 37602 32798
rect 36978 32734 36990 32786
rect 37042 32734 37054 32786
rect 33518 32722 33570 32734
rect 37550 32722 37602 32734
rect 38670 32786 38722 32798
rect 38670 32722 38722 32734
rect 39118 32786 39170 32798
rect 39118 32722 39170 32734
rect 39230 32786 39282 32798
rect 42254 32786 42306 32798
rect 39890 32734 39902 32786
rect 39954 32734 39966 32786
rect 39230 32722 39282 32734
rect 42254 32722 42306 32734
rect 42590 32786 42642 32798
rect 42590 32722 42642 32734
rect 43710 32786 43762 32798
rect 43710 32722 43762 32734
rect 44494 32786 44546 32798
rect 44494 32722 44546 32734
rect 45054 32786 45106 32798
rect 45054 32722 45106 32734
rect 49310 32786 49362 32798
rect 49310 32722 49362 32734
rect 49534 32786 49586 32798
rect 49858 32734 49870 32786
rect 49922 32783 49934 32786
rect 50082 32783 50094 32786
rect 49922 32737 50094 32783
rect 49922 32734 49934 32737
rect 50082 32734 50094 32737
rect 50146 32734 50158 32786
rect 49534 32722 49586 32734
rect 5742 32674 5794 32686
rect 5742 32610 5794 32622
rect 14926 32674 14978 32686
rect 14926 32610 14978 32622
rect 15150 32674 15202 32686
rect 15150 32610 15202 32622
rect 15486 32674 15538 32686
rect 15486 32610 15538 32622
rect 21870 32674 21922 32686
rect 21870 32610 21922 32622
rect 25790 32674 25842 32686
rect 25790 32610 25842 32622
rect 33406 32674 33458 32686
rect 33406 32610 33458 32622
rect 42478 32674 42530 32686
rect 52434 32622 52446 32674
rect 52498 32622 52510 32674
rect 42478 32610 42530 32622
rect 5630 32562 5682 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 5630 32498 5682 32510
rect 5966 32562 6018 32574
rect 21982 32562 22034 32574
rect 8754 32510 8766 32562
rect 8818 32510 8830 32562
rect 15922 32510 15934 32562
rect 15986 32510 15998 32562
rect 5966 32498 6018 32510
rect 21982 32498 22034 32510
rect 25454 32562 25506 32574
rect 25454 32498 25506 32510
rect 25902 32562 25954 32574
rect 25902 32498 25954 32510
rect 26238 32562 26290 32574
rect 26238 32498 26290 32510
rect 26574 32562 26626 32574
rect 26574 32498 26626 32510
rect 33742 32562 33794 32574
rect 37662 32562 37714 32574
rect 33954 32510 33966 32562
rect 34018 32510 34030 32562
rect 33742 32498 33794 32510
rect 37662 32498 37714 32510
rect 37774 32562 37826 32574
rect 37774 32498 37826 32510
rect 37886 32562 37938 32574
rect 39342 32562 39394 32574
rect 41806 32562 41858 32574
rect 38098 32510 38110 32562
rect 38162 32510 38174 32562
rect 38882 32510 38894 32562
rect 38946 32510 38958 32562
rect 39554 32510 39566 32562
rect 39618 32510 39630 32562
rect 40114 32510 40126 32562
rect 40178 32510 40190 32562
rect 37886 32498 37938 32510
rect 39342 32498 39394 32510
rect 41806 32498 41858 32510
rect 42030 32562 42082 32574
rect 42030 32498 42082 32510
rect 43598 32562 43650 32574
rect 43598 32498 43650 32510
rect 43934 32562 43986 32574
rect 43934 32498 43986 32510
rect 44158 32562 44210 32574
rect 44158 32498 44210 32510
rect 44942 32562 44994 32574
rect 44942 32498 44994 32510
rect 45614 32562 45666 32574
rect 53106 32510 53118 32562
rect 53170 32510 53182 32562
rect 45614 32498 45666 32510
rect 5182 32450 5234 32462
rect 15038 32450 15090 32462
rect 27022 32450 27074 32462
rect 43262 32450 43314 32462
rect 2482 32398 2494 32450
rect 2546 32398 2558 32450
rect 4610 32398 4622 32450
rect 4674 32398 4686 32450
rect 6402 32398 6414 32450
rect 6466 32398 6478 32450
rect 16258 32398 16270 32450
rect 16322 32398 16334 32450
rect 34738 32398 34750 32450
rect 34802 32398 34814 32450
rect 5182 32386 5234 32398
rect 15038 32386 15090 32398
rect 27022 32386 27074 32398
rect 43262 32386 43314 32398
rect 49086 32450 49138 32462
rect 49086 32386 49138 32398
rect 49422 32450 49474 32462
rect 50306 32398 50318 32450
rect 50370 32398 50382 32450
rect 49422 32386 49474 32398
rect 45054 32338 45106 32350
rect 45054 32274 45106 32286
rect 48862 32338 48914 32350
rect 49746 32286 49758 32338
rect 49810 32335 49822 32338
rect 50082 32335 50094 32338
rect 49810 32289 50094 32335
rect 49810 32286 49822 32289
rect 50082 32286 50094 32289
rect 50146 32286 50158 32338
rect 48862 32274 48914 32286
rect 1344 32170 53648 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 53648 32170
rect 1344 32084 53648 32118
rect 15150 32002 15202 32014
rect 15150 31938 15202 31950
rect 31726 32002 31778 32014
rect 50206 32002 50258 32014
rect 37202 31950 37214 32002
rect 37266 31999 37278 32002
rect 37538 31999 37550 32002
rect 37266 31953 37550 31999
rect 37266 31950 37278 31953
rect 37538 31950 37550 31953
rect 37602 31950 37614 32002
rect 31726 31938 31778 31950
rect 50206 31938 50258 31950
rect 5854 31890 5906 31902
rect 4946 31838 4958 31890
rect 5010 31838 5022 31890
rect 5854 31826 5906 31838
rect 7870 31890 7922 31902
rect 7870 31826 7922 31838
rect 9438 31890 9490 31902
rect 14478 31890 14530 31902
rect 37662 31890 37714 31902
rect 12674 31838 12686 31890
rect 12738 31838 12750 31890
rect 13682 31838 13694 31890
rect 13746 31838 13758 31890
rect 24994 31838 25006 31890
rect 25058 31838 25070 31890
rect 28466 31838 28478 31890
rect 28530 31838 28542 31890
rect 31042 31838 31054 31890
rect 31106 31838 31118 31890
rect 9438 31826 9490 31838
rect 14478 31826 14530 31838
rect 37662 31826 37714 31838
rect 38446 31890 38498 31902
rect 48514 31838 48526 31890
rect 48578 31838 48590 31890
rect 50530 31838 50542 31890
rect 50594 31838 50606 31890
rect 38446 31826 38498 31838
rect 5966 31778 6018 31790
rect 5058 31726 5070 31778
rect 5122 31726 5134 31778
rect 5966 31714 6018 31726
rect 6302 31778 6354 31790
rect 6302 31714 6354 31726
rect 7982 31778 8034 31790
rect 26350 31778 26402 31790
rect 9762 31726 9774 31778
rect 9826 31726 9838 31778
rect 13794 31726 13806 31778
rect 13858 31726 13870 31778
rect 15026 31726 15038 31778
rect 15090 31726 15102 31778
rect 16706 31726 16718 31778
rect 16770 31726 16782 31778
rect 23650 31726 23662 31778
rect 23714 31726 23726 31778
rect 24882 31726 24894 31778
rect 24946 31726 24958 31778
rect 7982 31714 8034 31726
rect 26350 31714 26402 31726
rect 26686 31778 26738 31790
rect 26686 31714 26738 31726
rect 26910 31778 26962 31790
rect 26910 31714 26962 31726
rect 27470 31778 27522 31790
rect 31390 31778 31442 31790
rect 27906 31726 27918 31778
rect 27970 31726 27982 31778
rect 28578 31726 28590 31778
rect 28642 31726 28654 31778
rect 27470 31714 27522 31726
rect 31390 31714 31442 31726
rect 32286 31778 32338 31790
rect 32286 31714 32338 31726
rect 33966 31778 34018 31790
rect 33966 31714 34018 31726
rect 34638 31778 34690 31790
rect 34638 31714 34690 31726
rect 39006 31778 39058 31790
rect 43374 31778 43426 31790
rect 39890 31726 39902 31778
rect 39954 31726 39966 31778
rect 45714 31726 45726 31778
rect 45778 31726 45790 31778
rect 39006 31714 39058 31726
rect 43374 31714 43426 31726
rect 4734 31666 4786 31678
rect 4734 31602 4786 31614
rect 5742 31666 5794 31678
rect 5742 31602 5794 31614
rect 6862 31666 6914 31678
rect 27358 31666 27410 31678
rect 10546 31614 10558 31666
rect 10610 31614 10622 31666
rect 15586 31614 15598 31666
rect 15650 31614 15662 31666
rect 16594 31614 16606 31666
rect 16658 31614 16670 31666
rect 24658 31614 24670 31666
rect 24722 31614 24734 31666
rect 6862 31602 6914 31614
rect 27358 31602 27410 31614
rect 31614 31666 31666 31678
rect 31614 31602 31666 31614
rect 31726 31666 31778 31678
rect 33394 31614 33406 31666
rect 33458 31614 33470 31666
rect 40562 31614 40574 31666
rect 40626 31614 40638 31666
rect 46386 31614 46398 31666
rect 46450 31614 46462 31666
rect 31726 31602 31778 31614
rect 6526 31554 6578 31566
rect 6526 31490 6578 31502
rect 6750 31554 6802 31566
rect 6750 31490 6802 31502
rect 7534 31554 7586 31566
rect 7534 31490 7586 31502
rect 7758 31554 7810 31566
rect 26014 31554 26066 31566
rect 23762 31502 23774 31554
rect 23826 31502 23838 31554
rect 7758 31490 7810 31502
rect 26014 31490 26066 31502
rect 26462 31554 26514 31566
rect 26462 31490 26514 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 28142 31554 28194 31566
rect 28142 31490 28194 31502
rect 28366 31554 28418 31566
rect 28366 31490 28418 31502
rect 29262 31554 29314 31566
rect 29262 31490 29314 31502
rect 30830 31554 30882 31566
rect 30830 31490 30882 31502
rect 31054 31554 31106 31566
rect 31054 31490 31106 31502
rect 33070 31554 33122 31566
rect 33070 31490 33122 31502
rect 34302 31554 34354 31566
rect 34302 31490 34354 31502
rect 34526 31554 34578 31566
rect 34526 31490 34578 31502
rect 37102 31554 37154 31566
rect 48974 31554 49026 31566
rect 42802 31502 42814 31554
rect 42866 31502 42878 31554
rect 37102 31490 37154 31502
rect 48974 31490 49026 31502
rect 49870 31554 49922 31566
rect 49870 31490 49922 31502
rect 50430 31554 50482 31566
rect 50430 31490 50482 31502
rect 1344 31386 53648 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 53648 31386
rect 1344 31300 53648 31334
rect 6638 31218 6690 31230
rect 6638 31154 6690 31166
rect 7534 31218 7586 31230
rect 7534 31154 7586 31166
rect 10110 31218 10162 31230
rect 10110 31154 10162 31166
rect 17726 31218 17778 31230
rect 26686 31218 26738 31230
rect 24322 31166 24334 31218
rect 24386 31166 24398 31218
rect 17726 31154 17778 31166
rect 26686 31154 26738 31166
rect 27358 31218 27410 31230
rect 31054 31218 31106 31230
rect 30482 31166 30494 31218
rect 30546 31166 30558 31218
rect 27358 31154 27410 31166
rect 31054 31154 31106 31166
rect 31278 31218 31330 31230
rect 31278 31154 31330 31166
rect 33966 31218 34018 31230
rect 33966 31154 34018 31166
rect 34526 31218 34578 31230
rect 34526 31154 34578 31166
rect 43822 31218 43874 31230
rect 43822 31154 43874 31166
rect 44382 31218 44434 31230
rect 44382 31154 44434 31166
rect 45278 31218 45330 31230
rect 45278 31154 45330 31166
rect 6078 31106 6130 31118
rect 6078 31042 6130 31054
rect 6190 31106 6242 31118
rect 21646 31106 21698 31118
rect 20402 31054 20414 31106
rect 20466 31054 20478 31106
rect 6190 31042 6242 31054
rect 21646 31042 21698 31054
rect 22094 31106 22146 31118
rect 22094 31042 22146 31054
rect 22542 31106 22594 31118
rect 22542 31042 22594 31054
rect 22654 31106 22706 31118
rect 22654 31042 22706 31054
rect 23438 31106 23490 31118
rect 27582 31106 27634 31118
rect 24210 31054 24222 31106
rect 24274 31054 24286 31106
rect 23438 31042 23490 31054
rect 27582 31042 27634 31054
rect 31838 31106 31890 31118
rect 31838 31042 31890 31054
rect 33630 31106 33682 31118
rect 33630 31042 33682 31054
rect 33742 31106 33794 31118
rect 33742 31042 33794 31054
rect 34302 31106 34354 31118
rect 34302 31042 34354 31054
rect 35310 31106 35362 31118
rect 35310 31042 35362 31054
rect 44830 31106 44882 31118
rect 44830 31042 44882 31054
rect 45054 31106 45106 31118
rect 52434 31054 52446 31106
rect 52498 31054 52510 31106
rect 45054 31042 45106 31054
rect 6526 30994 6578 31006
rect 6526 30930 6578 30942
rect 6750 30994 6802 31006
rect 6750 30930 6802 30942
rect 7198 30994 7250 31006
rect 7198 30930 7250 30942
rect 9774 30994 9826 31006
rect 9774 30930 9826 30942
rect 9998 30994 10050 31006
rect 9998 30930 10050 30942
rect 10222 30994 10274 31006
rect 21534 30994 21586 31006
rect 16034 30942 16046 30994
rect 16098 30942 16110 30994
rect 21074 30942 21086 30994
rect 21138 30942 21150 30994
rect 10222 30930 10274 30942
rect 21534 30930 21586 30942
rect 21758 30994 21810 31006
rect 21758 30930 21810 30942
rect 22318 30994 22370 31006
rect 27694 30994 27746 31006
rect 23538 30942 23550 30994
rect 23602 30942 23614 30994
rect 24098 30942 24110 30994
rect 24162 30942 24174 30994
rect 22318 30930 22370 30942
rect 27694 30930 27746 30942
rect 28142 30994 28194 31006
rect 28142 30930 28194 30942
rect 30830 30994 30882 31006
rect 30830 30930 30882 30942
rect 31390 30994 31442 31006
rect 31390 30930 31442 30942
rect 34190 30994 34242 31006
rect 34190 30930 34242 30942
rect 45390 30994 45442 31006
rect 53106 30942 53118 30994
rect 53170 30942 53182 30994
rect 45390 30930 45442 30942
rect 13134 30882 13186 30894
rect 16494 30882 16546 30894
rect 16370 30830 16382 30882
rect 16434 30830 16446 30882
rect 13134 30818 13186 30830
rect 16494 30818 16546 30830
rect 18286 30882 18338 30894
rect 18286 30818 18338 30830
rect 34862 30882 34914 30894
rect 34862 30818 34914 30830
rect 49982 30882 50034 30894
rect 50306 30830 50318 30882
rect 50370 30830 50382 30882
rect 49982 30818 50034 30830
rect 6078 30770 6130 30782
rect 7298 30718 7310 30770
rect 7362 30767 7374 30770
rect 7522 30767 7534 30770
rect 7362 30721 7534 30767
rect 7362 30718 7374 30721
rect 7522 30718 7534 30721
rect 7586 30718 7598 30770
rect 6078 30706 6130 30718
rect 1344 30602 53648 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 53648 30602
rect 1344 30516 53648 30550
rect 9886 30434 9938 30446
rect 9886 30370 9938 30382
rect 21982 30434 22034 30446
rect 21982 30370 22034 30382
rect 31278 30434 31330 30446
rect 31278 30370 31330 30382
rect 45166 30434 45218 30446
rect 45166 30370 45218 30382
rect 7198 30322 7250 30334
rect 28590 30322 28642 30334
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 15810 30270 15822 30322
rect 15874 30270 15886 30322
rect 17938 30270 17950 30322
rect 18002 30270 18014 30322
rect 24770 30270 24782 30322
rect 24834 30270 24846 30322
rect 43586 30270 43598 30322
rect 43650 30270 43662 30322
rect 7198 30258 7250 30270
rect 28590 30258 28642 30270
rect 5070 30210 5122 30222
rect 1698 30158 1710 30210
rect 1762 30158 1774 30210
rect 5070 30146 5122 30158
rect 6414 30210 6466 30222
rect 16158 30210 16210 30222
rect 9314 30158 9326 30210
rect 9378 30158 9390 30210
rect 15474 30158 15486 30210
rect 15538 30158 15550 30210
rect 6414 30146 6466 30158
rect 16158 30146 16210 30158
rect 16942 30210 16994 30222
rect 19406 30210 19458 30222
rect 18162 30158 18174 30210
rect 18226 30158 18238 30210
rect 16942 30146 16994 30158
rect 19406 30146 19458 30158
rect 22094 30210 22146 30222
rect 22094 30146 22146 30158
rect 22318 30210 22370 30222
rect 22318 30146 22370 30158
rect 22654 30210 22706 30222
rect 26126 30210 26178 30222
rect 23874 30158 23886 30210
rect 23938 30158 23950 30210
rect 24994 30158 25006 30210
rect 25058 30158 25070 30210
rect 22654 30146 22706 30158
rect 26126 30146 26178 30158
rect 29150 30210 29202 30222
rect 29150 30146 29202 30158
rect 31390 30210 31442 30222
rect 31390 30146 31442 30158
rect 42142 30210 42194 30222
rect 43374 30210 43426 30222
rect 43138 30158 43150 30210
rect 43202 30158 43214 30210
rect 42142 30146 42194 30158
rect 43374 30146 43426 30158
rect 6190 30098 6242 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 6190 30034 6242 30046
rect 6302 30098 6354 30110
rect 6302 30034 6354 30046
rect 6750 30098 6802 30110
rect 6750 30034 6802 30046
rect 17278 30098 17330 30110
rect 17278 30034 17330 30046
rect 18846 30098 18898 30110
rect 18846 30034 18898 30046
rect 22542 30098 22594 30110
rect 22542 30034 22594 30046
rect 23102 30098 23154 30110
rect 26462 30098 26514 30110
rect 24546 30046 24558 30098
rect 24610 30046 24622 30098
rect 25330 30046 25342 30098
rect 25394 30046 25406 30098
rect 23102 30034 23154 30046
rect 26462 30034 26514 30046
rect 29710 30098 29762 30110
rect 29710 30034 29762 30046
rect 45278 30098 45330 30110
rect 45278 30034 45330 30046
rect 52894 30098 52946 30110
rect 52894 30034 52946 30046
rect 53230 30098 53282 30110
rect 53230 30034 53282 30046
rect 9550 29986 9602 29998
rect 9550 29922 9602 29934
rect 9774 29986 9826 29998
rect 9774 29922 9826 29934
rect 21534 29986 21586 29998
rect 21534 29922 21586 29934
rect 21982 29986 22034 29998
rect 21982 29922 22034 29934
rect 23774 29986 23826 29998
rect 23774 29922 23826 29934
rect 25678 29986 25730 29998
rect 25678 29922 25730 29934
rect 26350 29986 26402 29998
rect 26350 29922 26402 29934
rect 27022 29986 27074 29998
rect 27022 29922 27074 29934
rect 28030 29986 28082 29998
rect 28030 29922 28082 29934
rect 30270 29986 30322 29998
rect 30270 29922 30322 29934
rect 31278 29986 31330 29998
rect 31278 29922 31330 29934
rect 31950 29986 32002 29998
rect 31950 29922 32002 29934
rect 39454 29986 39506 29998
rect 39454 29922 39506 29934
rect 40574 29986 40626 29998
rect 40574 29922 40626 29934
rect 42590 29986 42642 29998
rect 42590 29922 42642 29934
rect 43598 29986 43650 29998
rect 43598 29922 43650 29934
rect 43710 29986 43762 29998
rect 43710 29922 43762 29934
rect 45166 29986 45218 29998
rect 45166 29922 45218 29934
rect 45726 29986 45778 29998
rect 45726 29922 45778 29934
rect 1344 29818 53648 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 53648 29818
rect 1344 29732 53648 29766
rect 6862 29650 6914 29662
rect 6862 29586 6914 29598
rect 9998 29650 10050 29662
rect 9998 29586 10050 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 12910 29650 12962 29662
rect 31054 29650 31106 29662
rect 18946 29598 18958 29650
rect 19010 29598 19022 29650
rect 26898 29598 26910 29650
rect 26962 29598 26974 29650
rect 27906 29598 27918 29650
rect 27970 29598 27982 29650
rect 12910 29586 12962 29598
rect 31054 29586 31106 29598
rect 31502 29650 31554 29662
rect 31502 29586 31554 29598
rect 31726 29650 31778 29662
rect 35198 29650 35250 29662
rect 34178 29598 34190 29650
rect 34242 29598 34254 29650
rect 31726 29586 31778 29598
rect 35198 29586 35250 29598
rect 39230 29650 39282 29662
rect 39230 29586 39282 29598
rect 41134 29650 41186 29662
rect 41134 29586 41186 29598
rect 45502 29650 45554 29662
rect 45502 29586 45554 29598
rect 53342 29650 53394 29662
rect 53342 29586 53394 29598
rect 5854 29538 5906 29550
rect 5854 29474 5906 29486
rect 8654 29538 8706 29550
rect 8654 29474 8706 29486
rect 8878 29538 8930 29550
rect 8878 29474 8930 29486
rect 9662 29538 9714 29550
rect 18398 29538 18450 29550
rect 30718 29538 30770 29550
rect 11890 29486 11902 29538
rect 11954 29486 11966 29538
rect 18834 29486 18846 29538
rect 18898 29486 18910 29538
rect 20290 29486 20302 29538
rect 20354 29486 20366 29538
rect 27794 29486 27806 29538
rect 27858 29486 27870 29538
rect 9662 29474 9714 29486
rect 18398 29474 18450 29486
rect 30718 29474 30770 29486
rect 30830 29538 30882 29550
rect 30830 29474 30882 29486
rect 31278 29538 31330 29550
rect 31278 29474 31330 29486
rect 34526 29538 34578 29550
rect 34526 29474 34578 29486
rect 34974 29538 35026 29550
rect 34974 29474 35026 29486
rect 35534 29538 35586 29550
rect 35534 29474 35586 29486
rect 40126 29538 40178 29550
rect 40126 29474 40178 29486
rect 40350 29538 40402 29550
rect 47854 29538 47906 29550
rect 47394 29486 47406 29538
rect 47458 29486 47470 29538
rect 40350 29474 40402 29486
rect 47854 29474 47906 29486
rect 48190 29538 48242 29550
rect 51202 29486 51214 29538
rect 51266 29486 51278 29538
rect 48190 29474 48242 29486
rect 6414 29426 6466 29438
rect 6066 29374 6078 29426
rect 6130 29374 6142 29426
rect 6414 29362 6466 29374
rect 6750 29426 6802 29438
rect 6750 29362 6802 29374
rect 9886 29426 9938 29438
rect 9886 29362 9938 29374
rect 10446 29426 10498 29438
rect 10446 29362 10498 29374
rect 10782 29426 10834 29438
rect 10782 29362 10834 29374
rect 11006 29426 11058 29438
rect 18286 29426 18338 29438
rect 32174 29426 32226 29438
rect 12114 29374 12126 29426
rect 12178 29374 12190 29426
rect 13458 29374 13470 29426
rect 13522 29374 13534 29426
rect 17714 29374 17726 29426
rect 17778 29374 17790 29426
rect 18722 29374 18734 29426
rect 18786 29374 18798 29426
rect 20402 29374 20414 29426
rect 20466 29374 20478 29426
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 28242 29374 28254 29426
rect 28306 29374 28318 29426
rect 11006 29362 11058 29374
rect 18286 29362 18338 29374
rect 32174 29362 32226 29374
rect 34862 29426 34914 29438
rect 39678 29426 39730 29438
rect 35970 29374 35982 29426
rect 36034 29374 36046 29426
rect 34862 29362 34914 29374
rect 39678 29362 39730 29374
rect 40798 29426 40850 29438
rect 40798 29362 40850 29374
rect 41134 29426 41186 29438
rect 41134 29362 41186 29374
rect 41358 29426 41410 29438
rect 46510 29426 46562 29438
rect 42018 29374 42030 29426
rect 42082 29374 42094 29426
rect 41358 29362 41410 29374
rect 46510 29362 46562 29374
rect 46846 29426 46898 29438
rect 52446 29426 52498 29438
rect 51874 29374 51886 29426
rect 51938 29374 51950 29426
rect 46846 29362 46898 29374
rect 52446 29362 52498 29374
rect 6190 29314 6242 29326
rect 10894 29314 10946 29326
rect 8978 29262 8990 29314
rect 9042 29262 9054 29314
rect 6190 29250 6242 29262
rect 10894 29250 10946 29262
rect 12686 29314 12738 29326
rect 16830 29314 16882 29326
rect 13010 29262 13022 29314
rect 13074 29262 13086 29314
rect 14130 29262 14142 29314
rect 14194 29262 14206 29314
rect 16258 29262 16270 29314
rect 16322 29262 16334 29314
rect 12686 29250 12738 29262
rect 16830 29250 16882 29262
rect 26462 29314 26514 29326
rect 26462 29250 26514 29262
rect 28814 29314 28866 29326
rect 39902 29314 39954 29326
rect 44830 29314 44882 29326
rect 36642 29262 36654 29314
rect 36706 29262 36718 29314
rect 38770 29262 38782 29314
rect 38834 29262 38846 29314
rect 42690 29262 42702 29314
rect 42754 29262 42766 29314
rect 49074 29262 49086 29314
rect 49138 29262 49150 29314
rect 28814 29250 28866 29262
rect 39902 29250 39954 29262
rect 44830 29250 44882 29262
rect 6638 29202 6690 29214
rect 6638 29138 6690 29150
rect 31838 29202 31890 29214
rect 31838 29138 31890 29150
rect 47070 29202 47122 29214
rect 47070 29138 47122 29150
rect 1344 29034 53648 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 53648 29034
rect 1344 28948 53648 28982
rect 10110 28866 10162 28878
rect 40798 28866 40850 28878
rect 6402 28814 6414 28866
rect 6466 28814 6478 28866
rect 11778 28814 11790 28866
rect 11842 28814 11854 28866
rect 10110 28802 10162 28814
rect 40798 28802 40850 28814
rect 47070 28866 47122 28878
rect 47070 28802 47122 28814
rect 47406 28866 47458 28878
rect 47406 28802 47458 28814
rect 10222 28754 10274 28766
rect 10222 28690 10274 28702
rect 13694 28754 13746 28766
rect 13694 28690 13746 28702
rect 16494 28754 16546 28766
rect 16494 28690 16546 28702
rect 18286 28754 18338 28766
rect 18286 28690 18338 28702
rect 18734 28754 18786 28766
rect 18734 28690 18786 28702
rect 20302 28754 20354 28766
rect 20302 28690 20354 28702
rect 20750 28754 20802 28766
rect 20750 28690 20802 28702
rect 23214 28754 23266 28766
rect 23214 28690 23266 28702
rect 27022 28754 27074 28766
rect 34302 28754 34354 28766
rect 32162 28702 32174 28754
rect 32226 28702 32238 28754
rect 27022 28690 27074 28702
rect 34302 28690 34354 28702
rect 34974 28754 35026 28766
rect 34974 28690 35026 28702
rect 35870 28754 35922 28766
rect 35870 28690 35922 28702
rect 5742 28642 5794 28654
rect 8430 28642 8482 28654
rect 8194 28590 8206 28642
rect 8258 28590 8270 28642
rect 5742 28578 5794 28590
rect 8430 28578 8482 28590
rect 8542 28642 8594 28654
rect 8542 28578 8594 28590
rect 11454 28642 11506 28654
rect 18174 28642 18226 28654
rect 27582 28642 27634 28654
rect 36542 28642 36594 28654
rect 12002 28590 12014 28642
rect 12066 28590 12078 28642
rect 12898 28590 12910 28642
rect 12962 28590 12974 28642
rect 17602 28590 17614 28642
rect 17666 28590 17678 28642
rect 19618 28590 19630 28642
rect 19682 28590 19694 28642
rect 20066 28590 20078 28642
rect 20130 28590 20142 28642
rect 31378 28590 31390 28642
rect 31442 28590 31454 28642
rect 11454 28578 11506 28590
rect 18174 28578 18226 28590
rect 27582 28578 27634 28590
rect 36542 28578 36594 28590
rect 37214 28642 37266 28654
rect 37214 28578 37266 28590
rect 37438 28642 37490 28654
rect 37438 28578 37490 28590
rect 37550 28642 37602 28654
rect 37550 28578 37602 28590
rect 37774 28642 37826 28654
rect 37774 28578 37826 28590
rect 39678 28642 39730 28654
rect 39678 28578 39730 28590
rect 40462 28642 40514 28654
rect 40462 28578 40514 28590
rect 41358 28642 41410 28654
rect 48190 28642 48242 28654
rect 47954 28590 47966 28642
rect 48018 28590 48030 28642
rect 41358 28578 41410 28590
rect 48190 28578 48242 28590
rect 48302 28642 48354 28654
rect 48302 28578 48354 28590
rect 49086 28642 49138 28654
rect 49086 28578 49138 28590
rect 49646 28642 49698 28654
rect 49646 28578 49698 28590
rect 5854 28530 5906 28542
rect 5854 28466 5906 28478
rect 5966 28530 6018 28542
rect 22542 28530 22594 28542
rect 12786 28478 12798 28530
rect 12850 28478 12862 28530
rect 5966 28466 6018 28478
rect 22542 28466 22594 28478
rect 22654 28530 22706 28542
rect 22654 28466 22706 28478
rect 30942 28530 30994 28542
rect 30942 28466 30994 28478
rect 31054 28530 31106 28542
rect 31054 28466 31106 28478
rect 36206 28530 36258 28542
rect 36206 28466 36258 28478
rect 36318 28530 36370 28542
rect 36318 28466 36370 28478
rect 36990 28530 37042 28542
rect 36990 28466 37042 28478
rect 37998 28530 38050 28542
rect 37998 28466 38050 28478
rect 38110 28530 38162 28542
rect 38110 28466 38162 28478
rect 39342 28530 39394 28542
rect 39342 28466 39394 28478
rect 40126 28530 40178 28542
rect 40126 28466 40178 28478
rect 40686 28530 40738 28542
rect 40686 28466 40738 28478
rect 41806 28530 41858 28542
rect 46498 28478 46510 28530
rect 46562 28478 46574 28530
rect 46722 28478 46734 28530
rect 46786 28478 46798 28530
rect 41806 28466 41858 28478
rect 22878 28418 22930 28430
rect 8978 28366 8990 28418
rect 9042 28366 9054 28418
rect 22878 28354 22930 28366
rect 28030 28418 28082 28430
rect 28030 28354 28082 28366
rect 30494 28418 30546 28430
rect 30494 28354 30546 28366
rect 30718 28418 30770 28430
rect 30718 28354 30770 28366
rect 39006 28418 39058 28430
rect 39006 28354 39058 28366
rect 39454 28418 39506 28430
rect 39454 28354 39506 28366
rect 40238 28418 40290 28430
rect 40238 28354 40290 28366
rect 40798 28418 40850 28430
rect 48738 28366 48750 28418
rect 48802 28366 48814 28418
rect 40798 28354 40850 28366
rect 1344 28250 53648 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 53648 28250
rect 1344 28164 53648 28198
rect 6190 28082 6242 28094
rect 5966 28026 6018 28038
rect 5294 27970 5346 27982
rect 6190 28018 6242 28030
rect 7534 28082 7586 28094
rect 7534 28018 7586 28030
rect 8318 28082 8370 28094
rect 8318 28018 8370 28030
rect 21758 28082 21810 28094
rect 21758 28018 21810 28030
rect 22766 28082 22818 28094
rect 22766 28018 22818 28030
rect 23886 28082 23938 28094
rect 23886 28018 23938 28030
rect 24670 28082 24722 28094
rect 34526 28082 34578 28094
rect 34178 28030 34190 28082
rect 34242 28030 34254 28082
rect 24670 28018 24722 28030
rect 34526 28018 34578 28030
rect 34974 28082 35026 28094
rect 34974 28018 35026 28030
rect 35534 28082 35586 28094
rect 35534 28018 35586 28030
rect 35982 28082 36034 28094
rect 35982 28018 36034 28030
rect 36766 28082 36818 28094
rect 36766 28018 36818 28030
rect 40238 28082 40290 28094
rect 40238 28018 40290 28030
rect 40462 28082 40514 28094
rect 40462 28018 40514 28030
rect 41022 28082 41074 28094
rect 41022 28018 41074 28030
rect 45390 28082 45442 28094
rect 45390 28018 45442 28030
rect 46734 28082 46786 28094
rect 46734 28018 46786 28030
rect 47630 28082 47682 28094
rect 47630 28018 47682 28030
rect 48078 28082 48130 28094
rect 48078 28018 48130 28030
rect 48974 28082 49026 28094
rect 48974 28018 49026 28030
rect 5966 27962 6018 27974
rect 6638 27970 6690 27982
rect 5294 27906 5346 27918
rect 6638 27906 6690 27918
rect 7310 27970 7362 27982
rect 7310 27906 7362 27918
rect 7758 27970 7810 27982
rect 7758 27906 7810 27918
rect 10334 27970 10386 27982
rect 10334 27906 10386 27918
rect 10670 27970 10722 27982
rect 10670 27906 10722 27918
rect 19742 27970 19794 27982
rect 19742 27906 19794 27918
rect 21870 27970 21922 27982
rect 21870 27906 21922 27918
rect 23102 27970 23154 27982
rect 23102 27906 23154 27918
rect 23438 27970 23490 27982
rect 23438 27906 23490 27918
rect 24110 27970 24162 27982
rect 34862 27970 34914 27982
rect 31266 27918 31278 27970
rect 31330 27918 31342 27970
rect 24110 27906 24162 27918
rect 34862 27906 34914 27918
rect 45614 27970 45666 27982
rect 45614 27906 45666 27918
rect 46510 27970 46562 27982
rect 46510 27906 46562 27918
rect 4958 27858 5010 27870
rect 1698 27806 1710 27858
rect 1762 27806 1774 27858
rect 4958 27794 5010 27806
rect 5854 27858 5906 27870
rect 5854 27794 5906 27806
rect 6526 27858 6578 27870
rect 6526 27794 6578 27806
rect 6974 27858 7026 27870
rect 6974 27794 7026 27806
rect 7198 27858 7250 27870
rect 19630 27858 19682 27870
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 7198 27794 7250 27806
rect 19630 27794 19682 27806
rect 20190 27858 20242 27870
rect 20190 27794 20242 27806
rect 21534 27858 21586 27870
rect 21534 27794 21586 27806
rect 23550 27858 23602 27870
rect 23550 27794 23602 27806
rect 24222 27858 24274 27870
rect 40126 27858 40178 27870
rect 27234 27806 27246 27858
rect 27298 27806 27310 27858
rect 24222 27794 24274 27806
rect 40126 27794 40178 27806
rect 44270 27858 44322 27870
rect 45726 27858 45778 27870
rect 45042 27806 45054 27858
rect 45106 27806 45118 27858
rect 44270 27794 44322 27806
rect 45726 27794 45778 27806
rect 46398 27858 46450 27870
rect 53106 27806 53118 27858
rect 53170 27806 53182 27858
rect 46398 27794 46450 27806
rect 6862 27746 6914 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 6862 27682 6914 27694
rect 23214 27746 23266 27758
rect 23214 27682 23266 27694
rect 26910 27746 26962 27758
rect 26910 27682 26962 27694
rect 44606 27746 44658 27758
rect 44606 27682 44658 27694
rect 49982 27746 50034 27758
rect 50306 27694 50318 27746
rect 50370 27694 50382 27746
rect 52434 27694 52446 27746
rect 52498 27694 52510 27746
rect 49982 27682 50034 27694
rect 34974 27634 35026 27646
rect 34974 27570 35026 27582
rect 1344 27466 53648 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 53648 27466
rect 1344 27380 53648 27414
rect 6638 27298 6690 27310
rect 6638 27234 6690 27246
rect 27582 27298 27634 27310
rect 27582 27234 27634 27246
rect 37102 27298 37154 27310
rect 37102 27234 37154 27246
rect 45054 27298 45106 27310
rect 47518 27298 47570 27310
rect 45378 27246 45390 27298
rect 45442 27246 45454 27298
rect 45714 27246 45726 27298
rect 45778 27295 45790 27298
rect 46386 27295 46398 27298
rect 45778 27249 46398 27295
rect 45778 27246 45790 27249
rect 46386 27246 46398 27249
rect 46450 27246 46462 27298
rect 45054 27234 45106 27246
rect 47518 27234 47570 27246
rect 4846 27186 4898 27198
rect 4846 27122 4898 27134
rect 6526 27186 6578 27198
rect 16830 27186 16882 27198
rect 26014 27186 26066 27198
rect 16370 27134 16382 27186
rect 16434 27134 16446 27186
rect 23874 27134 23886 27186
rect 23938 27134 23950 27186
rect 6526 27122 6578 27134
rect 16830 27122 16882 27134
rect 26014 27122 26066 27134
rect 32286 27186 32338 27198
rect 32286 27122 32338 27134
rect 32734 27186 32786 27198
rect 32734 27122 32786 27134
rect 45950 27186 46002 27198
rect 45950 27122 46002 27134
rect 47630 27186 47682 27198
rect 47630 27122 47682 27134
rect 11006 27074 11058 27086
rect 11006 27010 11058 27022
rect 11342 27074 11394 27086
rect 11342 27010 11394 27022
rect 11678 27074 11730 27086
rect 21422 27074 21474 27086
rect 12226 27022 12238 27074
rect 12290 27022 12302 27074
rect 12450 27022 12462 27074
rect 12514 27022 12526 27074
rect 13458 27022 13470 27074
rect 13522 27022 13534 27074
rect 11678 27010 11730 27022
rect 21422 27010 21474 27022
rect 21646 27074 21698 27086
rect 21646 27010 21698 27022
rect 21982 27074 22034 27086
rect 30494 27074 30546 27086
rect 31838 27074 31890 27086
rect 23090 27022 23102 27074
rect 23154 27022 23166 27074
rect 31266 27022 31278 27074
rect 31330 27022 31342 27074
rect 21982 27010 22034 27022
rect 30494 27010 30546 27022
rect 31838 27010 31890 27022
rect 34526 27074 34578 27086
rect 36318 27074 36370 27086
rect 35074 27022 35086 27074
rect 35138 27022 35150 27074
rect 35634 27022 35646 27074
rect 35698 27022 35710 27074
rect 34526 27010 34578 27022
rect 36318 27010 36370 27022
rect 37214 27074 37266 27086
rect 40238 27074 40290 27086
rect 38434 27022 38446 27074
rect 38498 27022 38510 27074
rect 39106 27022 39118 27074
rect 39170 27022 39182 27074
rect 37214 27010 37266 27022
rect 40238 27010 40290 27022
rect 40686 27074 40738 27086
rect 40686 27010 40738 27022
rect 41470 27074 41522 27086
rect 41470 27010 41522 27022
rect 44830 27074 44882 27086
rect 44830 27010 44882 27022
rect 46622 27074 46674 27086
rect 53230 27074 53282 27086
rect 47058 27022 47070 27074
rect 47122 27022 47134 27074
rect 46622 27010 46674 27022
rect 53230 27010 53282 27022
rect 22206 26962 22258 26974
rect 14242 26910 14254 26962
rect 14306 26910 14318 26962
rect 22206 26898 22258 26910
rect 22542 26962 22594 26974
rect 22542 26898 22594 26910
rect 27694 26962 27746 26974
rect 27694 26898 27746 26910
rect 30606 26962 30658 26974
rect 30606 26898 30658 26910
rect 30718 26962 30770 26974
rect 30718 26898 30770 26910
rect 30830 26962 30882 26974
rect 30830 26898 30882 26910
rect 31726 26962 31778 26974
rect 37662 26962 37714 26974
rect 34850 26910 34862 26962
rect 34914 26910 34926 26962
rect 35858 26910 35870 26962
rect 35922 26910 35934 26962
rect 31726 26898 31778 26910
rect 37662 26898 37714 26910
rect 37998 26962 38050 26974
rect 40014 26962 40066 26974
rect 38658 26910 38670 26962
rect 38722 26910 38734 26962
rect 39330 26910 39342 26962
rect 39394 26910 39406 26962
rect 37998 26898 38050 26910
rect 40014 26898 40066 26910
rect 41022 26962 41074 26974
rect 41022 26898 41074 26910
rect 44270 26962 44322 26974
rect 44270 26898 44322 26910
rect 52894 26962 52946 26974
rect 52894 26898 52946 26910
rect 11230 26850 11282 26862
rect 11230 26786 11282 26798
rect 11902 26850 11954 26862
rect 11902 26786 11954 26798
rect 12014 26850 12066 26862
rect 12014 26786 12066 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 22430 26850 22482 26862
rect 22430 26786 22482 26798
rect 27582 26850 27634 26862
rect 27582 26786 27634 26798
rect 28142 26850 28194 26862
rect 28142 26786 28194 26798
rect 31502 26850 31554 26862
rect 31502 26786 31554 26798
rect 37102 26850 37154 26862
rect 37102 26786 37154 26798
rect 37886 26850 37938 26862
rect 37886 26786 37938 26798
rect 40126 26850 40178 26862
rect 40126 26786 40178 26798
rect 48078 26850 48130 26862
rect 48078 26786 48130 26798
rect 1344 26682 53648 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 53648 26682
rect 1344 26596 53648 26630
rect 6638 26514 6690 26526
rect 11678 26514 11730 26526
rect 9538 26462 9550 26514
rect 9602 26462 9614 26514
rect 6638 26450 6690 26462
rect 11678 26450 11730 26462
rect 15598 26514 15650 26526
rect 30942 26514 30994 26526
rect 24098 26462 24110 26514
rect 24162 26462 24174 26514
rect 26786 26462 26798 26514
rect 26850 26462 26862 26514
rect 15598 26450 15650 26462
rect 30942 26450 30994 26462
rect 49198 26514 49250 26526
rect 49198 26450 49250 26462
rect 51662 26514 51714 26526
rect 51662 26450 51714 26462
rect 53342 26514 53394 26526
rect 53342 26450 53394 26462
rect 5742 26402 5794 26414
rect 5742 26338 5794 26350
rect 6078 26402 6130 26414
rect 6078 26338 6130 26350
rect 12910 26402 12962 26414
rect 31166 26402 31218 26414
rect 15250 26350 15262 26402
rect 15314 26350 15326 26402
rect 29026 26350 29038 26402
rect 29090 26350 29102 26402
rect 12910 26338 12962 26350
rect 31166 26338 31218 26350
rect 45166 26402 45218 26414
rect 45166 26338 45218 26350
rect 49870 26402 49922 26414
rect 49870 26338 49922 26350
rect 6526 26290 6578 26302
rect 6526 26226 6578 26238
rect 6750 26290 6802 26302
rect 6750 26226 6802 26238
rect 7198 26290 7250 26302
rect 11566 26290 11618 26302
rect 9762 26238 9774 26290
rect 9826 26238 9838 26290
rect 11330 26238 11342 26290
rect 11394 26238 11406 26290
rect 7198 26226 7250 26238
rect 11566 26226 11618 26238
rect 11790 26290 11842 26302
rect 11790 26226 11842 26238
rect 11902 26290 11954 26302
rect 12574 26290 12626 26302
rect 18286 26290 18338 26302
rect 12338 26238 12350 26290
rect 12402 26238 12414 26290
rect 17714 26238 17726 26290
rect 17778 26238 17790 26290
rect 11902 26226 11954 26238
rect 12574 26226 12626 26238
rect 18286 26226 18338 26238
rect 24446 26290 24498 26302
rect 37774 26290 37826 26302
rect 29810 26238 29822 26290
rect 29874 26238 29886 26290
rect 31378 26238 31390 26290
rect 31442 26238 31454 26290
rect 31602 26238 31614 26290
rect 31666 26238 31678 26290
rect 24446 26226 24498 26238
rect 37774 26226 37826 26238
rect 39678 26290 39730 26302
rect 39678 26226 39730 26238
rect 40126 26290 40178 26302
rect 40126 26226 40178 26238
rect 40238 26290 40290 26302
rect 44606 26290 44658 26302
rect 43810 26238 43822 26290
rect 43874 26238 43886 26290
rect 40238 26226 40290 26238
rect 44606 26226 44658 26238
rect 49086 26290 49138 26302
rect 49086 26226 49138 26238
rect 49758 26290 49810 26302
rect 49758 26226 49810 26238
rect 51214 26290 51266 26302
rect 51874 26238 51886 26290
rect 51938 26238 51950 26290
rect 51214 26226 51266 26238
rect 13358 26178 13410 26190
rect 13358 26114 13410 26126
rect 18398 26178 18450 26190
rect 18398 26114 18450 26126
rect 18846 26178 18898 26190
rect 18846 26114 18898 26126
rect 22766 26178 22818 26190
rect 22766 26114 22818 26126
rect 30270 26178 30322 26190
rect 32174 26178 32226 26190
rect 31714 26126 31726 26178
rect 31778 26126 31790 26178
rect 30270 26114 30322 26126
rect 32174 26114 32226 26126
rect 39902 26178 39954 26190
rect 44270 26178 44322 26190
rect 40898 26126 40910 26178
rect 40962 26126 40974 26178
rect 43026 26126 43038 26178
rect 43090 26126 43102 26178
rect 39902 26114 39954 26126
rect 44270 26114 44322 26126
rect 12798 26066 12850 26078
rect 37998 26066 38050 26078
rect 49198 26066 49250 26078
rect 13122 26014 13134 26066
rect 13186 26063 13198 26066
rect 13346 26063 13358 26066
rect 13186 26017 13358 26063
rect 13186 26014 13198 26017
rect 13346 26014 13358 26017
rect 13410 26014 13422 26066
rect 38322 26014 38334 26066
rect 38386 26014 38398 26066
rect 12798 26002 12850 26014
rect 37998 26002 38050 26014
rect 49198 26002 49250 26014
rect 49870 26066 49922 26078
rect 49870 26002 49922 26014
rect 51550 26066 51602 26078
rect 51550 26002 51602 26014
rect 1344 25898 53648 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 53648 25898
rect 1344 25812 53648 25846
rect 6974 25730 7026 25742
rect 6974 25666 7026 25678
rect 19294 25730 19346 25742
rect 19294 25666 19346 25678
rect 19630 25730 19682 25742
rect 34850 25678 34862 25730
rect 34914 25727 34926 25730
rect 35186 25727 35198 25730
rect 34914 25681 35198 25727
rect 34914 25678 34926 25681
rect 35186 25678 35198 25681
rect 35250 25678 35262 25730
rect 19630 25666 19682 25678
rect 35198 25618 35250 25630
rect 6626 25566 6638 25618
rect 6690 25566 6702 25618
rect 31938 25566 31950 25618
rect 32002 25566 32014 25618
rect 34178 25566 34190 25618
rect 34242 25566 34254 25618
rect 35198 25554 35250 25566
rect 5854 25506 5906 25518
rect 5618 25454 5630 25506
rect 5682 25454 5694 25506
rect 5854 25442 5906 25454
rect 6078 25506 6130 25518
rect 8990 25506 9042 25518
rect 18622 25506 18674 25518
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 18386 25454 18398 25506
rect 18450 25454 18462 25506
rect 6078 25442 6130 25454
rect 8990 25442 9042 25454
rect 18622 25442 18674 25454
rect 19070 25506 19122 25518
rect 19070 25442 19122 25454
rect 19518 25506 19570 25518
rect 19518 25442 19570 25454
rect 25902 25506 25954 25518
rect 27694 25506 27746 25518
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 25902 25442 25954 25454
rect 27694 25442 27746 25454
rect 27918 25506 27970 25518
rect 27918 25442 27970 25454
rect 28142 25506 28194 25518
rect 49198 25506 49250 25518
rect 29362 25454 29374 25506
rect 29426 25454 29438 25506
rect 31266 25454 31278 25506
rect 31330 25454 31342 25506
rect 28142 25442 28194 25454
rect 49198 25442 49250 25454
rect 49870 25506 49922 25518
rect 49870 25442 49922 25454
rect 50878 25506 50930 25518
rect 50878 25442 50930 25454
rect 51102 25506 51154 25518
rect 51102 25442 51154 25454
rect 51662 25506 51714 25518
rect 51662 25442 51714 25454
rect 6750 25394 6802 25406
rect 10334 25394 10386 25406
rect 9426 25342 9438 25394
rect 9490 25342 9502 25394
rect 9650 25342 9662 25394
rect 9714 25342 9726 25394
rect 6750 25330 6802 25342
rect 10334 25330 10386 25342
rect 10670 25394 10722 25406
rect 10670 25330 10722 25342
rect 18958 25394 19010 25406
rect 26910 25394 26962 25406
rect 29934 25394 29986 25406
rect 26226 25342 26238 25394
rect 26290 25342 26302 25394
rect 29138 25342 29150 25394
rect 29202 25342 29214 25394
rect 18958 25330 19010 25342
rect 26910 25330 26962 25342
rect 29934 25330 29986 25342
rect 49646 25394 49698 25406
rect 49646 25330 49698 25342
rect 50206 25394 50258 25406
rect 50206 25330 50258 25342
rect 50430 25394 50482 25406
rect 50430 25330 50482 25342
rect 51326 25394 51378 25406
rect 51326 25330 51378 25342
rect 53230 25394 53282 25406
rect 53230 25330 53282 25342
rect 5966 25282 6018 25294
rect 25566 25282 25618 25294
rect 8978 25230 8990 25282
rect 9042 25230 9054 25282
rect 5966 25218 6018 25230
rect 25566 25218 25618 25230
rect 26798 25282 26850 25294
rect 30382 25282 30434 25294
rect 28466 25230 28478 25282
rect 28530 25230 28542 25282
rect 26798 25218 26850 25230
rect 30382 25218 30434 25230
rect 34750 25282 34802 25294
rect 34750 25218 34802 25230
rect 43374 25282 43426 25294
rect 43374 25218 43426 25230
rect 48414 25282 48466 25294
rect 48414 25218 48466 25230
rect 49534 25282 49586 25294
rect 49534 25218 49586 25230
rect 50542 25282 50594 25294
rect 50542 25218 50594 25230
rect 51550 25282 51602 25294
rect 51550 25218 51602 25230
rect 52894 25282 52946 25294
rect 52894 25218 52946 25230
rect 1344 25114 53648 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 53648 25114
rect 1344 25028 53648 25062
rect 5070 24946 5122 24958
rect 11454 24946 11506 24958
rect 5954 24894 5966 24946
rect 6018 24894 6030 24946
rect 6962 24894 6974 24946
rect 7026 24894 7038 24946
rect 5070 24882 5122 24894
rect 11454 24882 11506 24894
rect 13134 24946 13186 24958
rect 13134 24882 13186 24894
rect 18510 24946 18562 24958
rect 18510 24882 18562 24894
rect 19070 24946 19122 24958
rect 19070 24882 19122 24894
rect 29150 24946 29202 24958
rect 29150 24882 29202 24894
rect 30270 24946 30322 24958
rect 30270 24882 30322 24894
rect 34974 24946 35026 24958
rect 49086 24946 49138 24958
rect 42466 24894 42478 24946
rect 42530 24894 42542 24946
rect 43698 24894 43710 24946
rect 43762 24894 43774 24946
rect 34974 24882 35026 24894
rect 49086 24882 49138 24894
rect 50654 24946 50706 24958
rect 50654 24882 50706 24894
rect 51550 24946 51602 24958
rect 51550 24882 51602 24894
rect 11678 24834 11730 24846
rect 11678 24770 11730 24782
rect 12350 24834 12402 24846
rect 12350 24770 12402 24782
rect 13582 24834 13634 24846
rect 13582 24770 13634 24782
rect 18622 24834 18674 24846
rect 26126 24834 26178 24846
rect 22306 24782 22318 24834
rect 22370 24782 22382 24834
rect 18622 24770 18674 24782
rect 26126 24770 26178 24782
rect 28366 24834 28418 24846
rect 29710 24834 29762 24846
rect 34750 24834 34802 24846
rect 28578 24782 28590 24834
rect 28642 24782 28654 24834
rect 34402 24782 34414 24834
rect 34466 24782 34478 24834
rect 28366 24770 28418 24782
rect 29710 24770 29762 24782
rect 34750 24770 34802 24782
rect 48862 24834 48914 24846
rect 48862 24770 48914 24782
rect 50878 24834 50930 24846
rect 50878 24770 50930 24782
rect 5406 24722 5458 24734
rect 1698 24670 1710 24722
rect 1762 24670 1774 24722
rect 5406 24658 5458 24670
rect 5630 24722 5682 24734
rect 5630 24658 5682 24670
rect 6638 24722 6690 24734
rect 6638 24658 6690 24670
rect 11342 24722 11394 24734
rect 11342 24658 11394 24670
rect 11790 24722 11842 24734
rect 11790 24658 11842 24670
rect 12686 24722 12738 24734
rect 13470 24722 13522 24734
rect 13122 24670 13134 24722
rect 13186 24670 13198 24722
rect 12686 24658 12738 24670
rect 13470 24658 13522 24670
rect 18286 24722 18338 24734
rect 26462 24722 26514 24734
rect 29598 24722 29650 24734
rect 22978 24670 22990 24722
rect 23042 24670 23054 24722
rect 26898 24670 26910 24722
rect 26962 24670 26974 24722
rect 29026 24670 29038 24722
rect 29090 24670 29102 24722
rect 18286 24658 18338 24670
rect 26462 24658 26514 24670
rect 29598 24658 29650 24670
rect 30718 24722 30770 24734
rect 40350 24722 40402 24734
rect 42926 24722 42978 24734
rect 48750 24722 48802 24734
rect 34514 24670 34526 24722
rect 34578 24670 34590 24722
rect 35522 24670 35534 24722
rect 35586 24670 35598 24722
rect 38994 24670 39006 24722
rect 39058 24670 39070 24722
rect 42690 24670 42702 24722
rect 42754 24670 42766 24722
rect 45378 24670 45390 24722
rect 45442 24670 45454 24722
rect 30718 24658 30770 24670
rect 40350 24658 40402 24670
rect 42926 24658 42978 24670
rect 48750 24658 48802 24670
rect 49422 24722 49474 24734
rect 49422 24658 49474 24670
rect 50542 24722 50594 24734
rect 50542 24658 50594 24670
rect 51438 24722 51490 24734
rect 51438 24658 51490 24670
rect 51662 24722 51714 24734
rect 51662 24658 51714 24670
rect 51886 24722 51938 24734
rect 51886 24658 51938 24670
rect 53230 24722 53282 24734
rect 53230 24658 53282 24670
rect 12798 24610 12850 24622
rect 23662 24610 23714 24622
rect 2482 24558 2494 24610
rect 2546 24558 2558 24610
rect 4610 24558 4622 24610
rect 4674 24558 4686 24610
rect 11666 24558 11678 24610
rect 11730 24558 11742 24610
rect 20066 24558 20078 24610
rect 20130 24558 20142 24610
rect 12798 24546 12850 24558
rect 23662 24546 23714 24558
rect 26238 24610 26290 24622
rect 26238 24546 26290 24558
rect 27470 24610 27522 24622
rect 27470 24546 27522 24558
rect 28142 24610 28194 24622
rect 38334 24610 38386 24622
rect 39790 24610 39842 24622
rect 44270 24610 44322 24622
rect 34626 24558 34638 24610
rect 34690 24558 34702 24610
rect 36194 24558 36206 24610
rect 36258 24558 36270 24610
rect 39330 24558 39342 24610
rect 39394 24558 39406 24610
rect 42354 24558 42366 24610
rect 42418 24558 42430 24610
rect 28142 24546 28194 24558
rect 38334 24546 38386 24558
rect 39790 24546 39842 24558
rect 44270 24546 44322 24558
rect 44830 24610 44882 24622
rect 50206 24610 50258 24622
rect 46050 24558 46062 24610
rect 46114 24558 46126 24610
rect 48178 24558 48190 24610
rect 48242 24558 48254 24610
rect 44830 24546 44882 24558
rect 50206 24546 50258 24558
rect 29486 24498 29538 24510
rect 26674 24446 26686 24498
rect 26738 24446 26750 24498
rect 28914 24446 28926 24498
rect 28978 24446 28990 24498
rect 29486 24434 29538 24446
rect 44046 24498 44098 24510
rect 44046 24434 44098 24446
rect 1344 24330 53648 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 53648 24330
rect 1344 24244 53648 24278
rect 2606 24162 2658 24174
rect 2606 24098 2658 24110
rect 2942 24162 2994 24174
rect 2942 24098 2994 24110
rect 46622 24162 46674 24174
rect 46622 24098 46674 24110
rect 46958 24162 47010 24174
rect 46958 24098 47010 24110
rect 17278 24050 17330 24062
rect 14690 23998 14702 24050
rect 14754 23998 14766 24050
rect 16818 23998 16830 24050
rect 16882 23998 16894 24050
rect 17278 23986 17330 23998
rect 19070 24050 19122 24062
rect 27134 24050 27186 24062
rect 32062 24050 32114 24062
rect 22530 23998 22542 24050
rect 22594 23998 22606 24050
rect 24770 23998 24782 24050
rect 24834 23998 24846 24050
rect 29922 23998 29934 24050
rect 29986 23998 29998 24050
rect 19070 23986 19122 23998
rect 27134 23986 27186 23998
rect 32062 23986 32114 23998
rect 36206 24050 36258 24062
rect 36206 23986 36258 23998
rect 38782 24050 38834 24062
rect 38782 23986 38834 23998
rect 40798 24050 40850 24062
rect 44942 24050 44994 24062
rect 43810 23998 43822 24050
rect 43874 23998 43886 24050
rect 40798 23986 40850 23998
rect 44942 23986 44994 23998
rect 49870 24050 49922 24062
rect 49870 23986 49922 23998
rect 18958 23938 19010 23950
rect 34638 23938 34690 23950
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 11778 23886 11790 23938
rect 11842 23886 11854 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 29250 23886 29262 23938
rect 29314 23886 29326 23938
rect 18958 23874 19010 23886
rect 34638 23874 34690 23886
rect 34974 23938 35026 23950
rect 36318 23938 36370 23950
rect 35634 23886 35646 23938
rect 35698 23886 35710 23938
rect 34974 23874 35026 23886
rect 36318 23874 36370 23886
rect 37214 23938 37266 23950
rect 37214 23874 37266 23886
rect 41358 23938 41410 23950
rect 41358 23874 41410 23886
rect 43038 23938 43090 23950
rect 43038 23874 43090 23886
rect 44270 23938 44322 23950
rect 44270 23874 44322 23886
rect 45278 23938 45330 23950
rect 45278 23874 45330 23886
rect 50430 23938 50482 23950
rect 50430 23874 50482 23886
rect 35982 23826 36034 23838
rect 5618 23774 5630 23826
rect 5682 23774 5694 23826
rect 11554 23774 11566 23826
rect 11618 23774 11630 23826
rect 35982 23762 36034 23774
rect 36094 23826 36146 23838
rect 36094 23762 36146 23774
rect 36878 23826 36930 23838
rect 36878 23762 36930 23774
rect 42142 23826 42194 23838
rect 42142 23762 42194 23774
rect 46286 23826 46338 23838
rect 46286 23762 46338 23774
rect 46734 23826 46786 23838
rect 46734 23762 46786 23774
rect 50318 23826 50370 23838
rect 50318 23762 50370 23774
rect 2718 23714 2770 23726
rect 2718 23650 2770 23662
rect 3502 23714 3554 23726
rect 3502 23650 3554 23662
rect 5966 23714 6018 23726
rect 26014 23714 26066 23726
rect 8082 23662 8094 23714
rect 8146 23662 8158 23714
rect 5966 23650 6018 23662
rect 26014 23650 26066 23662
rect 28590 23714 28642 23726
rect 28590 23650 28642 23662
rect 34862 23714 34914 23726
rect 34862 23650 34914 23662
rect 37102 23714 37154 23726
rect 48190 23714 48242 23726
rect 45602 23662 45614 23714
rect 45666 23662 45678 23714
rect 37102 23650 37154 23662
rect 48190 23650 48242 23662
rect 50094 23714 50146 23726
rect 50094 23650 50146 23662
rect 50878 23714 50930 23726
rect 50878 23650 50930 23662
rect 1344 23546 53648 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 53648 23546
rect 1344 23460 53648 23494
rect 11230 23378 11282 23390
rect 6402 23326 6414 23378
rect 6466 23326 6478 23378
rect 11230 23314 11282 23326
rect 11454 23378 11506 23390
rect 11454 23314 11506 23326
rect 31614 23378 31666 23390
rect 31614 23314 31666 23326
rect 36542 23378 36594 23390
rect 36542 23314 36594 23326
rect 37214 23378 37266 23390
rect 37214 23314 37266 23326
rect 37774 23378 37826 23390
rect 49310 23378 49362 23390
rect 41234 23326 41246 23378
rect 41298 23326 41310 23378
rect 43586 23326 43598 23378
rect 43650 23326 43662 23378
rect 37774 23314 37826 23326
rect 49310 23314 49362 23326
rect 49758 23378 49810 23390
rect 49758 23314 49810 23326
rect 4846 23266 4898 23278
rect 4846 23202 4898 23214
rect 5070 23266 5122 23278
rect 5070 23202 5122 23214
rect 10110 23266 10162 23278
rect 10110 23202 10162 23214
rect 12686 23266 12738 23278
rect 12686 23202 12738 23214
rect 20078 23266 20130 23278
rect 39454 23266 39506 23278
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 20078 23202 20130 23214
rect 39454 23202 39506 23214
rect 10446 23154 10498 23166
rect 6178 23102 6190 23154
rect 6242 23102 6254 23154
rect 10446 23090 10498 23102
rect 10670 23154 10722 23166
rect 10670 23090 10722 23102
rect 10894 23154 10946 23166
rect 19518 23154 19570 23166
rect 21198 23154 21250 23166
rect 13010 23102 13022 23154
rect 13074 23102 13086 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 10894 23090 10946 23102
rect 19518 23090 19570 23102
rect 21198 23090 21250 23102
rect 31502 23154 31554 23166
rect 31502 23090 31554 23102
rect 37102 23154 37154 23166
rect 44046 23154 44098 23166
rect 41234 23102 41246 23154
rect 41298 23102 41310 23154
rect 41570 23102 41582 23154
rect 41634 23102 41646 23154
rect 42018 23102 42030 23154
rect 42082 23102 42094 23154
rect 43922 23102 43934 23154
rect 43986 23102 43998 23154
rect 37102 23090 37154 23102
rect 44046 23090 44098 23102
rect 44942 23154 44994 23166
rect 44942 23090 44994 23102
rect 48750 23154 48802 23166
rect 48750 23090 48802 23102
rect 49646 23154 49698 23166
rect 53106 23102 53118 23154
rect 53170 23102 53182 23154
rect 49646 23090 49698 23102
rect 4622 23042 4674 23054
rect 4622 22978 4674 22990
rect 10558 23042 10610 23054
rect 10558 22978 10610 22990
rect 27358 23042 27410 23054
rect 42590 23042 42642 23054
rect 45390 23042 45442 23054
rect 39330 22990 39342 23042
rect 39394 22990 39406 23042
rect 43474 22990 43486 23042
rect 43538 22990 43550 23042
rect 27358 22978 27410 22990
rect 42590 22978 42642 22990
rect 45390 22978 45442 22990
rect 47966 23042 48018 23054
rect 50306 22990 50318 23042
rect 50370 22990 50382 23042
rect 52434 22990 52446 23042
rect 52498 22990 52510 23042
rect 47966 22978 48018 22990
rect 5182 22930 5234 22942
rect 5182 22866 5234 22878
rect 11566 22930 11618 22942
rect 11566 22866 11618 22878
rect 13022 22930 13074 22942
rect 13022 22866 13074 22878
rect 37214 22930 37266 22942
rect 37214 22866 37266 22878
rect 39678 22930 39730 22942
rect 39678 22866 39730 22878
rect 49758 22930 49810 22942
rect 49758 22866 49810 22878
rect 1344 22762 53648 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 53648 22762
rect 1344 22676 53648 22710
rect 8318 22594 8370 22606
rect 8318 22530 8370 22542
rect 8990 22594 9042 22606
rect 8990 22530 9042 22542
rect 9550 22594 9602 22606
rect 15934 22594 15986 22606
rect 10546 22542 10558 22594
rect 10610 22542 10622 22594
rect 9550 22530 9602 22542
rect 15934 22530 15986 22542
rect 5070 22482 5122 22494
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 5070 22418 5122 22430
rect 7086 22482 7138 22494
rect 13694 22482 13746 22494
rect 9314 22430 9326 22482
rect 9378 22430 9390 22482
rect 7086 22418 7138 22430
rect 13694 22418 13746 22430
rect 18286 22482 18338 22494
rect 29934 22482 29986 22494
rect 27122 22430 27134 22482
rect 27186 22430 27198 22482
rect 18286 22418 18338 22430
rect 29934 22418 29986 22430
rect 31502 22482 31554 22494
rect 34750 22482 34802 22494
rect 43038 22482 43090 22494
rect 52782 22482 52834 22494
rect 32610 22430 32622 22482
rect 32674 22430 32686 22482
rect 41794 22430 41806 22482
rect 41858 22430 41870 22482
rect 47730 22430 47742 22482
rect 47794 22430 47806 22482
rect 49186 22430 49198 22482
rect 49250 22430 49262 22482
rect 31502 22418 31554 22430
rect 34750 22418 34802 22430
rect 43038 22418 43090 22430
rect 52782 22418 52834 22430
rect 8766 22370 8818 22382
rect 1698 22318 1710 22370
rect 1762 22318 1774 22370
rect 8306 22318 8318 22370
rect 8370 22318 8382 22370
rect 8766 22306 8818 22318
rect 9438 22370 9490 22382
rect 13918 22370 13970 22382
rect 10210 22318 10222 22370
rect 10274 22318 10286 22370
rect 10770 22318 10782 22370
rect 10834 22318 10846 22370
rect 9438 22306 9490 22318
rect 13918 22306 13970 22318
rect 14030 22370 14082 22382
rect 14814 22370 14866 22382
rect 27358 22370 27410 22382
rect 14354 22318 14366 22370
rect 14418 22318 14430 22370
rect 24322 22318 24334 22370
rect 24386 22318 24398 22370
rect 14030 22306 14082 22318
rect 14814 22306 14866 22318
rect 27358 22306 27410 22318
rect 27694 22370 27746 22382
rect 27694 22306 27746 22318
rect 28030 22370 28082 22382
rect 51326 22370 51378 22382
rect 29474 22318 29486 22370
rect 29538 22318 29550 22370
rect 31826 22318 31838 22370
rect 31890 22318 31902 22370
rect 37986 22318 37998 22370
rect 38050 22318 38062 22370
rect 39106 22318 39118 22370
rect 39170 22318 39182 22370
rect 41122 22318 41134 22370
rect 41186 22318 41198 22370
rect 42466 22318 42478 22370
rect 42530 22318 42542 22370
rect 44818 22318 44830 22370
rect 44882 22318 44894 22370
rect 48066 22318 48078 22370
rect 48130 22318 48142 22370
rect 28030 22306 28082 22318
rect 51326 22306 51378 22318
rect 5854 22258 5906 22270
rect 2482 22206 2494 22258
rect 2546 22206 2558 22258
rect 5854 22194 5906 22206
rect 6302 22258 6354 22270
rect 6302 22194 6354 22206
rect 7422 22258 7474 22270
rect 7422 22194 7474 22206
rect 7534 22258 7586 22270
rect 7534 22194 7586 22206
rect 7758 22258 7810 22270
rect 7758 22194 7810 22206
rect 7982 22258 8034 22270
rect 7982 22194 8034 22206
rect 9998 22258 10050 22270
rect 9998 22194 10050 22206
rect 13470 22258 13522 22270
rect 13470 22194 13522 22206
rect 16046 22258 16098 22270
rect 16046 22194 16098 22206
rect 18958 22258 19010 22270
rect 27582 22258 27634 22270
rect 50990 22258 51042 22270
rect 24994 22206 25006 22258
rect 25058 22206 25070 22258
rect 37314 22206 37326 22258
rect 37378 22206 37390 22258
rect 40562 22206 40574 22258
rect 40626 22206 40638 22258
rect 42130 22206 42142 22258
rect 42194 22206 42206 22258
rect 45602 22206 45614 22258
rect 45666 22206 45678 22258
rect 18958 22194 19010 22206
rect 27582 22194 27634 22206
rect 50990 22194 51042 22206
rect 51438 22258 51490 22270
rect 51438 22194 51490 22206
rect 51550 22258 51602 22270
rect 51550 22194 51602 22206
rect 52670 22258 52722 22270
rect 52670 22194 52722 22206
rect 5742 22146 5794 22158
rect 5742 22082 5794 22094
rect 5966 22146 6018 22158
rect 5966 22082 6018 22094
rect 6078 22146 6130 22158
rect 6078 22082 6130 22094
rect 10782 22146 10834 22158
rect 17726 22146 17778 22158
rect 14018 22094 14030 22146
rect 14082 22094 14094 22146
rect 10782 22082 10834 22094
rect 17726 22082 17778 22094
rect 18622 22146 18674 22158
rect 18622 22082 18674 22094
rect 30382 22146 30434 22158
rect 30382 22082 30434 22094
rect 36430 22146 36482 22158
rect 36430 22082 36482 22094
rect 41582 22146 41634 22158
rect 41582 22082 41634 22094
rect 43598 22146 43650 22158
rect 43598 22082 43650 22094
rect 44046 22146 44098 22158
rect 44046 22082 44098 22094
rect 52110 22146 52162 22158
rect 52110 22082 52162 22094
rect 52894 22146 52946 22158
rect 52894 22082 52946 22094
rect 1344 21978 53648 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 53648 21978
rect 1344 21892 53648 21926
rect 5406 21810 5458 21822
rect 5406 21746 5458 21758
rect 5742 21810 5794 21822
rect 5742 21746 5794 21758
rect 9550 21810 9602 21822
rect 9550 21746 9602 21758
rect 16830 21810 16882 21822
rect 16830 21746 16882 21758
rect 23886 21810 23938 21822
rect 23886 21746 23938 21758
rect 26910 21810 26962 21822
rect 26910 21746 26962 21758
rect 27134 21810 27186 21822
rect 27134 21746 27186 21758
rect 27582 21810 27634 21822
rect 27582 21746 27634 21758
rect 49982 21810 50034 21822
rect 49982 21746 50034 21758
rect 2718 21698 2770 21710
rect 2718 21634 2770 21646
rect 2942 21698 2994 21710
rect 2942 21634 2994 21646
rect 5854 21698 5906 21710
rect 5854 21634 5906 21646
rect 7310 21698 7362 21710
rect 7310 21634 7362 21646
rect 7422 21698 7474 21710
rect 7422 21634 7474 21646
rect 9662 21698 9714 21710
rect 39790 21698 39842 21710
rect 14242 21646 14254 21698
rect 14306 21646 14318 21698
rect 35298 21646 35310 21698
rect 35362 21646 35374 21698
rect 9662 21634 9714 21646
rect 39790 21634 39842 21646
rect 42366 21698 42418 21710
rect 42366 21634 42418 21646
rect 50430 21698 50482 21710
rect 50430 21634 50482 21646
rect 52670 21698 52722 21710
rect 52670 21634 52722 21646
rect 52894 21698 52946 21710
rect 52894 21634 52946 21646
rect 53230 21698 53282 21710
rect 53230 21634 53282 21646
rect 5630 21586 5682 21598
rect 5630 21522 5682 21534
rect 6526 21586 6578 21598
rect 6526 21522 6578 21534
rect 6638 21586 6690 21598
rect 17726 21586 17778 21598
rect 23998 21586 24050 21598
rect 26798 21586 26850 21598
rect 44046 21586 44098 21598
rect 49758 21586 49810 21598
rect 7074 21534 7086 21586
rect 7138 21534 7150 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 20626 21534 20638 21586
rect 20690 21534 20702 21586
rect 24322 21534 24334 21586
rect 24386 21534 24398 21586
rect 34850 21534 34862 21586
rect 34914 21534 34926 21586
rect 37090 21534 37102 21586
rect 37154 21534 37166 21586
rect 37762 21534 37774 21586
rect 37826 21534 37838 21586
rect 38098 21534 38110 21586
rect 38162 21534 38174 21586
rect 38658 21534 38670 21586
rect 38722 21534 38734 21586
rect 40226 21534 40238 21586
rect 40290 21534 40302 21586
rect 41570 21534 41582 21586
rect 41634 21534 41646 21586
rect 41794 21534 41806 21586
rect 41858 21534 41870 21586
rect 42802 21534 42814 21586
rect 42866 21534 42878 21586
rect 43138 21534 43150 21586
rect 43202 21534 43214 21586
rect 44482 21534 44494 21586
rect 44546 21534 44558 21586
rect 6638 21522 6690 21534
rect 17726 21522 17778 21534
rect 23998 21522 24050 21534
rect 3390 21474 3442 21486
rect 2594 21422 2606 21474
rect 2658 21422 2670 21474
rect 3390 21410 3442 21422
rect 4846 21474 4898 21486
rect 4846 21410 4898 21422
rect 6302 21474 6354 21486
rect 18286 21474 18338 21486
rect 16370 21422 16382 21474
rect 16434 21422 16446 21474
rect 21298 21422 21310 21474
rect 21362 21422 21374 21474
rect 23426 21422 23438 21474
rect 23490 21422 23502 21474
rect 6302 21410 6354 21422
rect 18286 21410 18338 21422
rect 6190 21362 6242 21374
rect 6190 21298 6242 21310
rect 23886 21362 23938 21374
rect 24337 21359 24383 21534
rect 26798 21522 26850 21534
rect 44046 21522 44098 21534
rect 49758 21522 49810 21534
rect 50094 21586 50146 21598
rect 50094 21522 50146 21534
rect 24446 21474 24498 21486
rect 24446 21410 24498 21422
rect 30718 21474 30770 21486
rect 30718 21410 30770 21422
rect 34302 21474 34354 21486
rect 34302 21410 34354 21422
rect 36206 21474 36258 21486
rect 45054 21474 45106 21486
rect 41234 21422 41246 21474
rect 41298 21422 41310 21474
rect 42690 21422 42702 21474
rect 42754 21422 42766 21474
rect 36206 21410 36258 21422
rect 45054 21410 45106 21422
rect 47742 21474 47794 21486
rect 47742 21410 47794 21422
rect 24434 21359 24446 21362
rect 24337 21313 24446 21359
rect 24434 21310 24446 21313
rect 24498 21310 24510 21362
rect 41010 21310 41022 21362
rect 41074 21310 41086 21362
rect 23886 21298 23938 21310
rect 1344 21194 53648 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 53648 21194
rect 1344 21108 53648 21142
rect 6638 21026 6690 21038
rect 43698 20974 43710 21026
rect 43762 21023 43774 21026
rect 43922 21023 43934 21026
rect 43762 20977 43934 21023
rect 43762 20974 43774 20977
rect 43922 20974 43934 20977
rect 43986 20974 43998 21026
rect 6638 20962 6690 20974
rect 6526 20914 6578 20926
rect 29934 20914 29986 20926
rect 43598 20914 43650 20926
rect 10770 20862 10782 20914
rect 10834 20862 10846 20914
rect 12898 20862 12910 20914
rect 12962 20862 12974 20914
rect 32946 20862 32958 20914
rect 33010 20862 33022 20914
rect 42018 20862 42030 20914
rect 42082 20862 42094 20914
rect 6526 20850 6578 20862
rect 29934 20850 29986 20862
rect 43598 20850 43650 20862
rect 5630 20802 5682 20814
rect 5630 20738 5682 20750
rect 6190 20802 6242 20814
rect 23886 20802 23938 20814
rect 31166 20802 31218 20814
rect 34862 20802 34914 20814
rect 45166 20802 45218 20814
rect 9986 20750 9998 20802
rect 10050 20750 10062 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 30370 20750 30382 20802
rect 30434 20750 30446 20802
rect 31826 20750 31838 20802
rect 31890 20750 31902 20802
rect 33506 20750 33518 20802
rect 33570 20750 33582 20802
rect 37986 20750 37998 20802
rect 38050 20750 38062 20802
rect 39106 20750 39118 20802
rect 39170 20750 39182 20802
rect 41458 20750 41470 20802
rect 41522 20750 41534 20802
rect 42130 20750 42142 20802
rect 42194 20750 42206 20802
rect 42466 20750 42478 20802
rect 42530 20750 42542 20802
rect 44930 20750 44942 20802
rect 44994 20750 45006 20802
rect 6190 20738 6242 20750
rect 23886 20738 23938 20750
rect 31166 20738 31218 20750
rect 34862 20738 34914 20750
rect 45166 20738 45218 20750
rect 45390 20802 45442 20814
rect 45390 20738 45442 20750
rect 45950 20802 46002 20814
rect 45950 20738 46002 20750
rect 5966 20690 6018 20702
rect 5966 20626 6018 20638
rect 23214 20690 23266 20702
rect 23214 20626 23266 20638
rect 23438 20690 23490 20702
rect 23438 20626 23490 20638
rect 29150 20690 29202 20702
rect 29150 20626 29202 20638
rect 30830 20690 30882 20702
rect 32050 20638 32062 20690
rect 32114 20638 32126 20690
rect 37314 20638 37326 20690
rect 37378 20638 37390 20690
rect 40562 20638 40574 20690
rect 40626 20638 40638 20690
rect 30830 20626 30882 20638
rect 5742 20578 5794 20590
rect 5742 20514 5794 20526
rect 9662 20578 9714 20590
rect 23550 20578 23602 20590
rect 16594 20526 16606 20578
rect 16658 20526 16670 20578
rect 9662 20514 9714 20526
rect 23550 20514 23602 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 29486 20578 29538 20590
rect 29486 20514 29538 20526
rect 30942 20578 30994 20590
rect 41582 20578 41634 20590
rect 31490 20526 31502 20578
rect 31554 20526 31566 20578
rect 34514 20526 34526 20578
rect 34578 20526 34590 20578
rect 30942 20514 30994 20526
rect 41582 20514 41634 20526
rect 41694 20578 41746 20590
rect 41694 20514 41746 20526
rect 43934 20578 43986 20590
rect 43934 20514 43986 20526
rect 45054 20578 45106 20590
rect 45054 20514 45106 20526
rect 49534 20578 49586 20590
rect 50430 20578 50482 20590
rect 49858 20526 49870 20578
rect 49922 20526 49934 20578
rect 49534 20514 49586 20526
rect 50430 20514 50482 20526
rect 1344 20410 53648 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 53648 20410
rect 1344 20324 53648 20358
rect 5854 20242 5906 20254
rect 5854 20178 5906 20190
rect 41918 20242 41970 20254
rect 41918 20178 41970 20190
rect 42254 20242 42306 20254
rect 42254 20178 42306 20190
rect 47406 20242 47458 20254
rect 47406 20178 47458 20190
rect 2830 20130 2882 20142
rect 2830 20066 2882 20078
rect 3054 20130 3106 20142
rect 3054 20066 3106 20078
rect 3502 20130 3554 20142
rect 3502 20066 3554 20078
rect 7870 20130 7922 20142
rect 7870 20066 7922 20078
rect 8094 20130 8146 20142
rect 8094 20066 8146 20078
rect 9550 20130 9602 20142
rect 9550 20066 9602 20078
rect 14702 20130 14754 20142
rect 14702 20066 14754 20078
rect 15038 20130 15090 20142
rect 15710 20130 15762 20142
rect 15362 20078 15374 20130
rect 15426 20078 15438 20130
rect 15038 20066 15090 20078
rect 15710 20066 15762 20078
rect 16494 20130 16546 20142
rect 16494 20066 16546 20078
rect 16830 20130 16882 20142
rect 16830 20066 16882 20078
rect 23998 20130 24050 20142
rect 33182 20130 33234 20142
rect 26786 20078 26798 20130
rect 26850 20078 26862 20130
rect 30482 20078 30494 20130
rect 30546 20078 30558 20130
rect 31826 20078 31838 20130
rect 31890 20078 31902 20130
rect 23998 20066 24050 20078
rect 33182 20066 33234 20078
rect 37214 20130 37266 20142
rect 37214 20066 37266 20078
rect 37438 20130 37490 20142
rect 37438 20066 37490 20078
rect 40126 20130 40178 20142
rect 40126 20066 40178 20078
rect 41806 20130 41858 20142
rect 41806 20066 41858 20078
rect 42814 20130 42866 20142
rect 44606 20130 44658 20142
rect 44034 20078 44046 20130
rect 44098 20078 44110 20130
rect 42814 20066 42866 20078
rect 44606 20066 44658 20078
rect 44830 20130 44882 20142
rect 44830 20066 44882 20078
rect 45390 20130 45442 20142
rect 45390 20066 45442 20078
rect 45502 20130 45554 20142
rect 45502 20066 45554 20078
rect 46734 20130 46786 20142
rect 46734 20066 46786 20078
rect 46958 20130 47010 20142
rect 48862 20130 48914 20142
rect 47506 20078 47518 20130
rect 47570 20078 47582 20130
rect 49746 20078 49758 20130
rect 49810 20078 49822 20130
rect 46958 20066 47010 20078
rect 48862 20066 48914 20078
rect 5182 20018 5234 20030
rect 8206 20018 8258 20030
rect 5618 19966 5630 20018
rect 5682 19966 5694 20018
rect 5182 19954 5234 19966
rect 8206 19954 8258 19966
rect 9886 20018 9938 20030
rect 9886 19954 9938 19966
rect 10334 20018 10386 20030
rect 23774 20018 23826 20030
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 17490 19966 17502 20018
rect 17554 19966 17566 20018
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 10334 19954 10386 19966
rect 23774 19954 23826 19966
rect 24110 20018 24162 20030
rect 24110 19954 24162 19966
rect 26126 20018 26178 20030
rect 32174 20018 32226 20030
rect 26562 19966 26574 20018
rect 26626 19966 26638 20018
rect 30258 19966 30270 20018
rect 30322 19966 30334 20018
rect 26126 19954 26178 19966
rect 32174 19954 32226 19966
rect 32398 20018 32450 20030
rect 32398 19954 32450 19966
rect 37102 20018 37154 20030
rect 37102 19954 37154 19966
rect 39790 20018 39842 20030
rect 39790 19954 39842 19966
rect 40014 20018 40066 20030
rect 40014 19954 40066 19966
rect 41470 20018 41522 20030
rect 44494 20018 44546 20030
rect 43810 19966 43822 20018
rect 43874 19966 43886 20018
rect 41470 19954 41522 19966
rect 44494 19954 44546 19966
rect 44942 20018 44994 20030
rect 44942 19954 44994 19966
rect 45614 20018 45666 20030
rect 45614 19954 45666 19966
rect 46286 20018 46338 20030
rect 46286 19954 46338 19966
rect 47294 20018 47346 20030
rect 49422 20018 49474 20030
rect 48066 19966 48078 20018
rect 48130 19966 48142 20018
rect 50306 19966 50318 20018
rect 50370 19966 50382 20018
rect 47294 19954 47346 19966
rect 49422 19954 49474 19966
rect 8654 19906 8706 19918
rect 8654 19842 8706 19854
rect 11118 19906 11170 19918
rect 11118 19842 11170 19854
rect 16270 19906 16322 19918
rect 24558 19906 24610 19918
rect 18162 19854 18174 19906
rect 18226 19854 18238 19906
rect 20290 19854 20302 19906
rect 20354 19854 20366 19906
rect 21410 19854 21422 19906
rect 21474 19854 21486 19906
rect 23538 19854 23550 19906
rect 23602 19854 23614 19906
rect 16270 19842 16322 19854
rect 24558 19842 24610 19854
rect 30942 19906 30994 19918
rect 37886 19906 37938 19918
rect 42366 19906 42418 19918
rect 46062 19906 46114 19918
rect 33058 19854 33070 19906
rect 33122 19854 33134 19906
rect 41010 19854 41022 19906
rect 41074 19854 41086 19906
rect 43474 19854 43486 19906
rect 43538 19854 43550 19906
rect 30942 19842 30994 19854
rect 37886 19842 37938 19854
rect 42366 19842 42418 19854
rect 46062 19842 46114 19854
rect 46510 19906 46562 19918
rect 51090 19854 51102 19906
rect 51154 19854 51166 19906
rect 53218 19854 53230 19906
rect 53282 19854 53294 19906
rect 46510 19842 46562 19854
rect 2718 19794 2770 19806
rect 2718 19730 2770 19742
rect 10222 19794 10274 19806
rect 10222 19730 10274 19742
rect 33406 19794 33458 19806
rect 48750 19794 48802 19806
rect 37538 19742 37550 19794
rect 37602 19791 37614 19794
rect 37874 19791 37886 19794
rect 37602 19745 37886 19791
rect 37602 19742 37614 19745
rect 37874 19742 37886 19745
rect 37938 19742 37950 19794
rect 47842 19742 47854 19794
rect 47906 19742 47918 19794
rect 33406 19730 33458 19742
rect 48750 19730 48802 19742
rect 49086 19794 49138 19806
rect 49086 19730 49138 19742
rect 1344 19626 53648 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 53648 19626
rect 1344 19540 53648 19574
rect 8430 19458 8482 19470
rect 8430 19394 8482 19406
rect 8766 19458 8818 19470
rect 8766 19394 8818 19406
rect 5182 19346 5234 19358
rect 17054 19346 17106 19358
rect 2482 19294 2494 19346
rect 2546 19294 2558 19346
rect 4610 19294 4622 19346
rect 4674 19294 4686 19346
rect 11666 19294 11678 19346
rect 11730 19294 11742 19346
rect 5182 19282 5234 19294
rect 17054 19282 17106 19294
rect 23886 19346 23938 19358
rect 23886 19282 23938 19294
rect 32846 19346 32898 19358
rect 39230 19346 39282 19358
rect 37202 19294 37214 19346
rect 37266 19294 37278 19346
rect 32846 19282 32898 19294
rect 39230 19282 39282 19294
rect 47070 19346 47122 19358
rect 52222 19346 52274 19358
rect 49298 19294 49310 19346
rect 49362 19294 49374 19346
rect 47070 19282 47122 19294
rect 52222 19282 52274 19294
rect 20526 19234 20578 19246
rect 23774 19234 23826 19246
rect 1698 19182 1710 19234
rect 1762 19182 1774 19234
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 20526 19170 20578 19182
rect 23774 19170 23826 19182
rect 23998 19234 24050 19246
rect 29374 19234 29426 19246
rect 25442 19182 25454 19234
rect 25506 19182 25518 19234
rect 23998 19170 24050 19182
rect 29374 19170 29426 19182
rect 30270 19234 30322 19246
rect 30270 19170 30322 19182
rect 33630 19234 33682 19246
rect 41246 19234 41298 19246
rect 53230 19234 53282 19246
rect 37538 19182 37550 19234
rect 37602 19182 37614 19234
rect 41570 19182 41582 19234
rect 41634 19182 41646 19234
rect 48178 19182 48190 19234
rect 48242 19182 48254 19234
rect 33630 19170 33682 19182
rect 41246 19170 41298 19182
rect 53230 19170 53282 19182
rect 11454 19122 11506 19134
rect 11454 19058 11506 19070
rect 24334 19122 24386 19134
rect 37998 19122 38050 19134
rect 42142 19122 42194 19134
rect 26226 19070 26238 19122
rect 26290 19070 26302 19122
rect 39554 19070 39566 19122
rect 39618 19070 39630 19122
rect 47730 19070 47742 19122
rect 47794 19070 47806 19122
rect 24334 19058 24386 19070
rect 37998 19058 38050 19070
rect 42142 19058 42194 19070
rect 8654 19010 8706 19022
rect 23102 19010 23154 19022
rect 20178 18958 20190 19010
rect 20242 18958 20254 19010
rect 8654 18946 8706 18958
rect 23102 18946 23154 18958
rect 24782 19010 24834 19022
rect 29038 19010 29090 19022
rect 25106 18958 25118 19010
rect 25170 18958 25182 19010
rect 28466 18958 28478 19010
rect 28530 18958 28542 19010
rect 24782 18946 24834 18958
rect 29038 18946 29090 18958
rect 29262 19010 29314 19022
rect 29262 18946 29314 18958
rect 29822 19010 29874 19022
rect 29822 18946 29874 18958
rect 33742 19010 33794 19022
rect 33742 18946 33794 18958
rect 33966 19010 34018 19022
rect 33966 18946 34018 18958
rect 34302 19010 34354 19022
rect 34302 18946 34354 18958
rect 38782 19010 38834 19022
rect 43822 19010 43874 19022
rect 40562 18958 40574 19010
rect 40626 18958 40638 19010
rect 38782 18946 38834 18958
rect 43822 18946 43874 18958
rect 44270 19010 44322 19022
rect 44270 18946 44322 18958
rect 44942 19010 44994 19022
rect 44942 18946 44994 18958
rect 45390 19010 45442 19022
rect 45390 18946 45442 18958
rect 47406 19010 47458 19022
rect 47406 18946 47458 18958
rect 52894 19010 52946 19022
rect 52894 18946 52946 18958
rect 1344 18842 53648 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 53648 18842
rect 1344 18756 53648 18790
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 32398 18674 32450 18686
rect 32398 18610 32450 18622
rect 50990 18674 51042 18686
rect 50990 18610 51042 18622
rect 8766 18562 8818 18574
rect 6066 18510 6078 18562
rect 6130 18510 6142 18562
rect 7970 18510 7982 18562
rect 8034 18510 8046 18562
rect 8766 18498 8818 18510
rect 27134 18562 27186 18574
rect 31726 18562 31778 18574
rect 31378 18510 31390 18562
rect 31442 18510 31454 18562
rect 27134 18498 27186 18510
rect 31726 18498 31778 18510
rect 31950 18562 32002 18574
rect 31950 18498 32002 18510
rect 32510 18562 32562 18574
rect 32510 18498 32562 18510
rect 38110 18562 38162 18574
rect 38110 18498 38162 18510
rect 39118 18562 39170 18574
rect 41246 18562 41298 18574
rect 46622 18562 46674 18574
rect 51438 18562 51490 18574
rect 40114 18510 40126 18562
rect 40178 18510 40190 18562
rect 43810 18510 43822 18562
rect 43874 18510 43886 18562
rect 49634 18510 49646 18562
rect 49698 18510 49710 18562
rect 39118 18498 39170 18510
rect 41246 18498 41298 18510
rect 46622 18498 46674 18510
rect 51438 18498 51490 18510
rect 8318 18450 8370 18462
rect 6738 18398 6750 18450
rect 6802 18398 6814 18450
rect 7522 18398 7534 18450
rect 7586 18398 7598 18450
rect 8318 18386 8370 18398
rect 8990 18450 9042 18462
rect 16270 18450 16322 18462
rect 12562 18398 12574 18450
rect 12626 18398 12638 18450
rect 8990 18386 9042 18398
rect 16270 18386 16322 18398
rect 26910 18450 26962 18462
rect 26910 18386 26962 18398
rect 27022 18450 27074 18462
rect 27022 18386 27074 18398
rect 27582 18450 27634 18462
rect 32174 18450 32226 18462
rect 41470 18450 41522 18462
rect 31490 18398 31502 18450
rect 31554 18398 31566 18450
rect 33170 18398 33182 18450
rect 33234 18398 33246 18450
rect 37090 18398 37102 18450
rect 37154 18398 37166 18450
rect 38434 18398 38446 18450
rect 38498 18398 38510 18450
rect 38882 18398 38894 18450
rect 38946 18398 38958 18450
rect 39778 18398 39790 18450
rect 39842 18398 39854 18450
rect 27582 18386 27634 18398
rect 32174 18386 32226 18398
rect 41470 18386 41522 18398
rect 41694 18450 41746 18462
rect 41694 18386 41746 18398
rect 41918 18450 41970 18462
rect 41918 18386 41970 18398
rect 42590 18450 42642 18462
rect 42590 18386 42642 18398
rect 43150 18450 43202 18462
rect 43150 18386 43202 18398
rect 43486 18450 43538 18462
rect 43486 18386 43538 18398
rect 45166 18450 45218 18462
rect 51774 18450 51826 18462
rect 46946 18398 46958 18450
rect 47010 18398 47022 18450
rect 49410 18398 49422 18450
rect 49474 18398 49486 18450
rect 50754 18398 50766 18450
rect 50818 18398 50830 18450
rect 45166 18386 45218 18398
rect 51774 18386 51826 18398
rect 51886 18450 51938 18462
rect 51886 18386 51938 18398
rect 52222 18450 52274 18462
rect 52222 18386 52274 18398
rect 52446 18450 52498 18462
rect 52446 18386 52498 18398
rect 52558 18450 52610 18462
rect 52558 18386 52610 18398
rect 52894 18450 52946 18462
rect 52894 18386 52946 18398
rect 9662 18338 9714 18350
rect 15710 18338 15762 18350
rect 6626 18286 6638 18338
rect 6690 18286 6702 18338
rect 8642 18286 8654 18338
rect 8706 18286 8718 18338
rect 13234 18286 13246 18338
rect 13298 18286 13310 18338
rect 15362 18286 15374 18338
rect 15426 18286 15438 18338
rect 9662 18274 9714 18286
rect 15710 18274 15762 18286
rect 25342 18338 25394 18350
rect 25342 18274 25394 18286
rect 26574 18338 26626 18350
rect 35982 18338 36034 18350
rect 37774 18338 37826 18350
rect 44606 18338 44658 18350
rect 31602 18286 31614 18338
rect 31666 18286 31678 18338
rect 33842 18286 33854 18338
rect 33906 18286 33918 18338
rect 37426 18286 37438 18338
rect 37490 18286 37502 18338
rect 40226 18286 40238 18338
rect 40290 18286 40302 18338
rect 26574 18274 26626 18286
rect 35982 18274 36034 18286
rect 37774 18274 37826 18286
rect 44606 18274 44658 18286
rect 46734 18338 46786 18350
rect 46734 18274 46786 18286
rect 47854 18338 47906 18350
rect 47854 18274 47906 18286
rect 51550 18338 51602 18350
rect 51550 18274 51602 18286
rect 15822 18226 15874 18238
rect 15822 18162 15874 18174
rect 38446 18226 38498 18238
rect 38446 18162 38498 18174
rect 42366 18226 42418 18238
rect 42366 18162 42418 18174
rect 51102 18226 51154 18238
rect 51102 18162 51154 18174
rect 1344 18058 53648 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 53648 18058
rect 1344 17972 53648 18006
rect 9886 17890 9938 17902
rect 9886 17826 9938 17838
rect 32622 17890 32674 17902
rect 32622 17826 32674 17838
rect 42478 17890 42530 17902
rect 42478 17826 42530 17838
rect 51214 17890 51266 17902
rect 51214 17826 51266 17838
rect 9102 17778 9154 17790
rect 9102 17714 9154 17726
rect 10110 17778 10162 17790
rect 10110 17714 10162 17726
rect 10670 17778 10722 17790
rect 36542 17778 36594 17790
rect 20738 17726 20750 17778
rect 20802 17726 20814 17778
rect 29922 17726 29934 17778
rect 29986 17726 29998 17778
rect 33618 17726 33630 17778
rect 33682 17726 33694 17778
rect 40674 17726 40686 17778
rect 40738 17726 40750 17778
rect 43698 17726 43710 17778
rect 43762 17726 43774 17778
rect 46610 17726 46622 17778
rect 46674 17726 46686 17778
rect 48738 17726 48750 17778
rect 48802 17726 48814 17778
rect 10670 17714 10722 17726
rect 36542 17714 36594 17726
rect 5630 17666 5682 17678
rect 5630 17602 5682 17614
rect 5854 17666 5906 17678
rect 6862 17666 6914 17678
rect 6178 17614 6190 17666
rect 6242 17614 6254 17666
rect 5854 17602 5906 17614
rect 6862 17602 6914 17614
rect 7422 17666 7474 17678
rect 7422 17602 7474 17614
rect 8654 17666 8706 17678
rect 34414 17666 34466 17678
rect 49198 17666 49250 17678
rect 9650 17614 9662 17666
rect 9714 17614 9726 17666
rect 17826 17614 17838 17666
rect 17890 17614 17902 17666
rect 29138 17614 29150 17666
rect 29202 17614 29214 17666
rect 33954 17614 33966 17666
rect 34018 17614 34030 17666
rect 38994 17614 39006 17666
rect 39058 17614 39070 17666
rect 39554 17614 39566 17666
rect 39618 17614 39630 17666
rect 43138 17614 43150 17666
rect 43202 17614 43214 17666
rect 45938 17614 45950 17666
rect 46002 17614 46014 17666
rect 8654 17602 8706 17614
rect 34414 17602 34466 17614
rect 49198 17602 49250 17614
rect 51998 17666 52050 17678
rect 51998 17602 52050 17614
rect 6526 17554 6578 17566
rect 6526 17490 6578 17502
rect 10222 17554 10274 17566
rect 25790 17554 25842 17566
rect 18610 17502 18622 17554
rect 18674 17502 18686 17554
rect 10222 17490 10274 17502
rect 25790 17490 25842 17502
rect 32734 17554 32786 17566
rect 32734 17490 32786 17502
rect 33182 17554 33234 17566
rect 42590 17554 42642 17566
rect 33842 17502 33854 17554
rect 33906 17502 33918 17554
rect 39218 17502 39230 17554
rect 39282 17502 39294 17554
rect 33182 17490 33234 17502
rect 42590 17490 42642 17502
rect 44158 17554 44210 17566
rect 44158 17490 44210 17502
rect 50542 17554 50594 17566
rect 50542 17490 50594 17502
rect 50654 17554 50706 17566
rect 50654 17490 50706 17502
rect 51102 17554 51154 17566
rect 51102 17490 51154 17502
rect 51214 17554 51266 17566
rect 51214 17490 51266 17502
rect 51662 17554 51714 17566
rect 51662 17490 51714 17502
rect 51774 17554 51826 17566
rect 51774 17490 51826 17502
rect 6638 17442 6690 17454
rect 6638 17378 6690 17390
rect 7086 17442 7138 17454
rect 17054 17442 17106 17454
rect 8306 17390 8318 17442
rect 8370 17390 8382 17442
rect 7086 17378 7138 17390
rect 17054 17378 17106 17390
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 24894 17442 24946 17454
rect 24894 17378 24946 17390
rect 25454 17442 25506 17454
rect 25454 17378 25506 17390
rect 25678 17442 25730 17454
rect 25678 17378 25730 17390
rect 28590 17442 28642 17454
rect 34190 17442 34242 17454
rect 32162 17390 32174 17442
rect 32226 17390 32238 17442
rect 28590 17378 28642 17390
rect 34190 17378 34242 17390
rect 38110 17442 38162 17454
rect 38110 17378 38162 17390
rect 38558 17442 38610 17454
rect 44942 17442 44994 17454
rect 42914 17390 42926 17442
rect 42978 17390 42990 17442
rect 38558 17378 38610 17390
rect 44942 17378 44994 17390
rect 45502 17442 45554 17454
rect 45502 17378 45554 17390
rect 50878 17442 50930 17454
rect 50878 17378 50930 17390
rect 1344 17274 53648 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 53648 17274
rect 1344 17188 53648 17222
rect 6414 17106 6466 17118
rect 6414 17042 6466 17054
rect 7534 17106 7586 17118
rect 7534 17042 7586 17054
rect 13134 17106 13186 17118
rect 13134 17042 13186 17054
rect 15822 17106 15874 17118
rect 15822 17042 15874 17054
rect 18174 17106 18226 17118
rect 18174 17042 18226 17054
rect 24222 17106 24274 17118
rect 24222 17042 24274 17054
rect 32286 17106 32338 17118
rect 32286 17042 32338 17054
rect 36430 17106 36482 17118
rect 36430 17042 36482 17054
rect 37998 17106 38050 17118
rect 37998 17042 38050 17054
rect 51326 17106 51378 17118
rect 51326 17042 51378 17054
rect 51774 17106 51826 17118
rect 51774 17042 51826 17054
rect 13918 16994 13970 17006
rect 2482 16942 2494 16994
rect 2546 16942 2558 16994
rect 13918 16930 13970 16942
rect 14478 16994 14530 17006
rect 14478 16930 14530 16942
rect 17390 16994 17442 17006
rect 24334 16994 24386 17006
rect 40014 16994 40066 17006
rect 17602 16942 17614 16994
rect 17666 16942 17678 16994
rect 20290 16942 20302 16994
rect 20354 16991 20366 16994
rect 20626 16991 20638 16994
rect 20354 16945 20638 16991
rect 20354 16942 20366 16945
rect 20626 16942 20638 16945
rect 20690 16942 20702 16994
rect 39218 16942 39230 16994
rect 39282 16942 39294 16994
rect 17390 16930 17442 16942
rect 24334 16930 24386 16942
rect 40014 16930 40066 16942
rect 45054 16994 45106 17006
rect 45054 16930 45106 16942
rect 49310 16994 49362 17006
rect 49310 16930 49362 16942
rect 52894 16994 52946 17006
rect 52894 16930 52946 16942
rect 5070 16882 5122 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 5070 16818 5122 16830
rect 6302 16882 6354 16894
rect 13470 16882 13522 16894
rect 6514 16830 6526 16882
rect 6578 16830 6590 16882
rect 7074 16830 7086 16882
rect 7138 16830 7150 16882
rect 13122 16830 13134 16882
rect 13186 16830 13198 16882
rect 6302 16818 6354 16830
rect 13470 16818 13522 16830
rect 13582 16882 13634 16894
rect 13582 16818 13634 16830
rect 14590 16882 14642 16894
rect 14590 16818 14642 16830
rect 14814 16882 14866 16894
rect 16046 16882 16098 16894
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 14814 16818 14866 16830
rect 16046 16818 16098 16830
rect 16382 16882 16434 16894
rect 20078 16882 20130 16894
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 17938 16830 17950 16882
rect 18002 16830 18014 16882
rect 16382 16818 16434 16830
rect 20078 16818 20130 16830
rect 20190 16882 20242 16894
rect 23998 16882 24050 16894
rect 36318 16882 36370 16894
rect 20962 16830 20974 16882
rect 21026 16830 21038 16882
rect 25218 16830 25230 16882
rect 25282 16830 25294 16882
rect 20190 16818 20242 16830
rect 23998 16818 24050 16830
rect 36318 16818 36370 16830
rect 38558 16882 38610 16894
rect 44494 16882 44546 16894
rect 38770 16830 38782 16882
rect 38834 16830 38846 16882
rect 40226 16830 40238 16882
rect 40290 16830 40302 16882
rect 43138 16830 43150 16882
rect 43202 16830 43214 16882
rect 38558 16818 38610 16830
rect 44494 16818 44546 16830
rect 49198 16882 49250 16894
rect 49198 16818 49250 16830
rect 49534 16882 49586 16894
rect 49534 16818 49586 16830
rect 52670 16882 52722 16894
rect 52670 16818 52722 16830
rect 53230 16882 53282 16894
rect 53230 16818 53282 16830
rect 16158 16770 16210 16782
rect 4610 16718 4622 16770
rect 4674 16718 4686 16770
rect 16158 16706 16210 16718
rect 17838 16770 17890 16782
rect 21634 16718 21646 16770
rect 21698 16718 21710 16770
rect 23762 16718 23774 16770
rect 23826 16718 23838 16770
rect 26002 16718 26014 16770
rect 26066 16718 26078 16770
rect 28130 16718 28142 16770
rect 28194 16718 28206 16770
rect 39218 16718 39230 16770
rect 39282 16718 39294 16770
rect 42578 16718 42590 16770
rect 42642 16718 42654 16770
rect 17838 16706 17890 16718
rect 14926 16658 14978 16670
rect 6850 16606 6862 16658
rect 6914 16606 6926 16658
rect 14926 16594 14978 16606
rect 16494 16658 16546 16670
rect 16494 16594 16546 16606
rect 1344 16490 53648 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 53648 16490
rect 1344 16404 53648 16438
rect 15374 16322 15426 16334
rect 44706 16270 44718 16322
rect 44770 16319 44782 16322
rect 44930 16319 44942 16322
rect 44770 16273 44942 16319
rect 44770 16270 44782 16273
rect 44930 16270 44942 16273
rect 44994 16270 45006 16322
rect 15374 16258 15426 16270
rect 12798 16210 12850 16222
rect 6066 16158 6078 16210
rect 6130 16158 6142 16210
rect 12450 16158 12462 16210
rect 12514 16158 12526 16210
rect 12798 16146 12850 16158
rect 17390 16210 17442 16222
rect 44270 16210 44322 16222
rect 34850 16158 34862 16210
rect 34914 16158 34926 16210
rect 42018 16158 42030 16210
rect 42082 16158 42094 16210
rect 17390 16146 17442 16158
rect 44270 16146 44322 16158
rect 44942 16210 44994 16222
rect 44942 16146 44994 16158
rect 51214 16210 51266 16222
rect 51214 16146 51266 16158
rect 4958 16098 5010 16110
rect 6862 16098 6914 16110
rect 13582 16098 13634 16110
rect 4610 16046 4622 16098
rect 4674 16046 4686 16098
rect 6178 16046 6190 16098
rect 6242 16046 6254 16098
rect 9650 16046 9662 16098
rect 9714 16046 9726 16098
rect 4958 16034 5010 16046
rect 6862 16034 6914 16046
rect 13582 16034 13634 16046
rect 15710 16098 15762 16110
rect 15710 16034 15762 16046
rect 23102 16098 23154 16110
rect 23102 16034 23154 16046
rect 23662 16098 23714 16110
rect 25118 16098 25170 16110
rect 24434 16046 24446 16098
rect 24498 16046 24510 16098
rect 23662 16034 23714 16046
rect 25118 16034 25170 16046
rect 25678 16098 25730 16110
rect 48638 16098 48690 16110
rect 34962 16046 34974 16098
rect 35026 16046 35038 16098
rect 37538 16046 37550 16098
rect 37602 16046 37614 16098
rect 38994 16046 39006 16098
rect 39058 16046 39070 16098
rect 39442 16046 39454 16098
rect 39506 16046 39518 16098
rect 40226 16046 40238 16098
rect 40290 16046 40302 16098
rect 41234 16046 41246 16098
rect 41298 16046 41310 16098
rect 42354 16046 42366 16098
rect 42418 16046 42430 16098
rect 43810 16046 43822 16098
rect 43874 16046 43886 16098
rect 25678 16034 25730 16046
rect 48638 16034 48690 16046
rect 48862 16098 48914 16110
rect 48862 16034 48914 16046
rect 49534 16098 49586 16110
rect 49534 16034 49586 16046
rect 50094 16098 50146 16110
rect 50094 16034 50146 16046
rect 50766 16098 50818 16110
rect 50766 16034 50818 16046
rect 51886 16098 51938 16110
rect 51886 16034 51938 16046
rect 52222 16098 52274 16110
rect 52222 16034 52274 16046
rect 52894 16098 52946 16110
rect 52894 16034 52946 16046
rect 53118 16098 53170 16110
rect 53118 16034 53170 16046
rect 5070 15986 5122 15998
rect 5070 15922 5122 15934
rect 6526 15986 6578 15998
rect 6526 15922 6578 15934
rect 6638 15986 6690 15998
rect 15486 15986 15538 15998
rect 10322 15934 10334 15986
rect 10386 15934 10398 15986
rect 6638 15922 6690 15934
rect 15486 15922 15538 15934
rect 17278 15986 17330 15998
rect 17278 15922 17330 15934
rect 17502 15986 17554 15998
rect 17502 15922 17554 15934
rect 23214 15986 23266 15998
rect 23214 15922 23266 15934
rect 24670 15986 24722 15998
rect 24670 15922 24722 15934
rect 25342 15986 25394 15998
rect 25342 15922 25394 15934
rect 35646 15986 35698 15998
rect 49198 15986 49250 15998
rect 38546 15934 38558 15986
rect 38610 15934 38622 15986
rect 35646 15922 35698 15934
rect 49198 15922 49250 15934
rect 49758 15986 49810 15998
rect 49758 15922 49810 15934
rect 49982 15986 50034 15998
rect 49982 15922 50034 15934
rect 50430 15986 50482 15998
rect 50430 15922 50482 15934
rect 52670 15986 52722 15998
rect 52670 15922 52722 15934
rect 12910 15874 12962 15886
rect 12910 15810 12962 15822
rect 23326 15874 23378 15886
rect 23326 15810 23378 15822
rect 23998 15874 24050 15886
rect 23998 15810 24050 15822
rect 25566 15874 25618 15886
rect 48750 15874 48802 15886
rect 37650 15822 37662 15874
rect 37714 15822 37726 15874
rect 38434 15822 38446 15874
rect 38498 15822 38510 15874
rect 25566 15810 25618 15822
rect 48750 15810 48802 15822
rect 50654 15874 50706 15886
rect 50654 15810 50706 15822
rect 51998 15874 52050 15886
rect 51998 15810 52050 15822
rect 52782 15874 52834 15886
rect 52782 15810 52834 15822
rect 1344 15706 53648 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 53648 15706
rect 1344 15620 53648 15654
rect 6302 15538 6354 15550
rect 6302 15474 6354 15486
rect 10446 15538 10498 15550
rect 10446 15474 10498 15486
rect 18174 15538 18226 15550
rect 35310 15538 35362 15550
rect 40238 15538 40290 15550
rect 28802 15486 28814 15538
rect 28866 15486 28878 15538
rect 34290 15486 34302 15538
rect 34354 15486 34366 15538
rect 39218 15486 39230 15538
rect 39282 15486 39294 15538
rect 18174 15474 18226 15486
rect 35310 15474 35362 15486
rect 40238 15474 40290 15486
rect 41022 15538 41074 15550
rect 52334 15538 52386 15550
rect 45490 15486 45502 15538
rect 45554 15486 45566 15538
rect 46498 15486 46510 15538
rect 46562 15486 46574 15538
rect 41022 15474 41074 15486
rect 52334 15474 52386 15486
rect 5966 15426 6018 15438
rect 5966 15362 6018 15374
rect 6078 15426 6130 15438
rect 10334 15426 10386 15438
rect 13582 15426 13634 15438
rect 8642 15374 8654 15426
rect 8706 15374 8718 15426
rect 10546 15374 10558 15426
rect 10610 15374 10622 15426
rect 6078 15362 6130 15374
rect 10334 15362 10386 15374
rect 13582 15362 13634 15374
rect 13918 15426 13970 15438
rect 13918 15362 13970 15374
rect 14254 15426 14306 15438
rect 14254 15362 14306 15374
rect 14590 15426 14642 15438
rect 14590 15362 14642 15374
rect 17390 15426 17442 15438
rect 33406 15426 33458 15438
rect 17602 15374 17614 15426
rect 17666 15374 17678 15426
rect 19506 15374 19518 15426
rect 19570 15374 19582 15426
rect 17390 15362 17442 15374
rect 33406 15362 33458 15374
rect 33966 15426 34018 15438
rect 48750 15426 48802 15438
rect 36418 15374 36430 15426
rect 36482 15374 36494 15426
rect 38770 15374 38782 15426
rect 38834 15374 38846 15426
rect 33966 15362 34018 15374
rect 48750 15362 48802 15374
rect 51774 15426 51826 15438
rect 51774 15362 51826 15374
rect 22094 15314 22146 15326
rect 8418 15262 8430 15314
rect 8482 15262 8494 15314
rect 11106 15262 11118 15314
rect 11170 15262 11182 15314
rect 17938 15262 17950 15314
rect 18002 15262 18014 15314
rect 18834 15262 18846 15314
rect 18898 15262 18910 15314
rect 22094 15250 22146 15262
rect 28478 15314 28530 15326
rect 28478 15250 28530 15262
rect 29150 15314 29202 15326
rect 44718 15314 44770 15326
rect 29586 15262 29598 15314
rect 29650 15262 29662 15314
rect 36082 15262 36094 15314
rect 36146 15262 36158 15314
rect 37314 15262 37326 15314
rect 37378 15262 37390 15314
rect 39330 15262 39342 15314
rect 39394 15262 39406 15314
rect 44146 15262 44158 15314
rect 44210 15262 44222 15314
rect 29150 15250 29202 15262
rect 44718 15250 44770 15262
rect 45838 15314 45890 15326
rect 51102 15314 51154 15326
rect 46274 15262 46286 15314
rect 46338 15262 46350 15314
rect 49074 15262 49086 15314
rect 49138 15262 49150 15314
rect 45838 15250 45890 15262
rect 51102 15250 51154 15262
rect 51438 15314 51490 15326
rect 51438 15250 51490 15262
rect 33518 15202 33570 15214
rect 48862 15202 48914 15214
rect 21634 15150 21646 15202
rect 21698 15150 21710 15202
rect 30370 15150 30382 15202
rect 30434 15150 30446 15202
rect 32498 15150 32510 15202
rect 32562 15150 32574 15202
rect 41346 15150 41358 15202
rect 41410 15150 41422 15202
rect 43474 15150 43486 15202
rect 43538 15150 43550 15202
rect 33518 15138 33570 15150
rect 48862 15138 48914 15150
rect 51326 15202 51378 15214
rect 51326 15138 51378 15150
rect 52110 15202 52162 15214
rect 52110 15138 52162 15150
rect 52222 15202 52274 15214
rect 52222 15138 52274 15150
rect 17838 15090 17890 15102
rect 10882 15038 10894 15090
rect 10946 15038 10958 15090
rect 17838 15026 17890 15038
rect 1344 14922 53648 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 53648 14922
rect 1344 14836 53648 14870
rect 6414 14754 6466 14766
rect 6414 14690 6466 14702
rect 6638 14754 6690 14766
rect 6638 14690 6690 14702
rect 36094 14754 36146 14766
rect 36094 14690 36146 14702
rect 42254 14754 42306 14766
rect 42254 14690 42306 14702
rect 9662 14642 9714 14654
rect 9662 14578 9714 14590
rect 29374 14642 29426 14654
rect 29374 14578 29426 14590
rect 31166 14642 31218 14654
rect 42702 14642 42754 14654
rect 40786 14590 40798 14642
rect 40850 14590 40862 14642
rect 31166 14578 31218 14590
rect 42702 14578 42754 14590
rect 45838 14642 45890 14654
rect 52670 14642 52722 14654
rect 48850 14590 48862 14642
rect 48914 14590 48926 14642
rect 50978 14590 50990 14642
rect 51042 14590 51054 14642
rect 45838 14578 45890 14590
rect 52670 14578 52722 14590
rect 8094 14530 8146 14542
rect 6178 14478 6190 14530
rect 6242 14478 6254 14530
rect 8094 14466 8146 14478
rect 8318 14530 8370 14542
rect 8878 14530 8930 14542
rect 8642 14478 8654 14530
rect 8706 14478 8718 14530
rect 8318 14466 8370 14478
rect 8878 14466 8930 14478
rect 9214 14530 9266 14542
rect 15710 14530 15762 14542
rect 17614 14530 17666 14542
rect 19070 14530 19122 14542
rect 15138 14478 15150 14530
rect 15202 14478 15214 14530
rect 17378 14478 17390 14530
rect 17442 14478 17454 14530
rect 17714 14478 17726 14530
rect 17778 14478 17790 14530
rect 9214 14466 9266 14478
rect 15710 14466 15762 14478
rect 17614 14466 17666 14478
rect 19070 14466 19122 14478
rect 24334 14530 24386 14542
rect 24334 14466 24386 14478
rect 26014 14530 26066 14542
rect 31838 14530 31890 14542
rect 31490 14478 31502 14530
rect 31554 14478 31566 14530
rect 32050 14478 32062 14530
rect 32114 14478 32126 14530
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 42242 14478 42254 14530
rect 42306 14478 42318 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 46274 14478 46286 14530
rect 46338 14478 46350 14530
rect 48178 14478 48190 14530
rect 48242 14478 48254 14530
rect 26014 14466 26066 14478
rect 31838 14466 31890 14478
rect 6750 14418 6802 14430
rect 17166 14418 17218 14430
rect 15362 14366 15374 14418
rect 15426 14366 15438 14418
rect 6750 14354 6802 14366
rect 17166 14354 17218 14366
rect 18286 14418 18338 14430
rect 18286 14354 18338 14366
rect 18398 14418 18450 14430
rect 18398 14354 18450 14366
rect 32286 14418 32338 14430
rect 32286 14354 32338 14366
rect 35982 14418 36034 14430
rect 41918 14418 41970 14430
rect 38770 14366 38782 14418
rect 38834 14366 38846 14418
rect 39666 14366 39678 14418
rect 39730 14366 39742 14418
rect 35982 14354 36034 14366
rect 41918 14354 41970 14366
rect 46958 14418 47010 14430
rect 46958 14354 47010 14366
rect 8206 14306 8258 14318
rect 8206 14242 8258 14254
rect 9102 14306 9154 14318
rect 9102 14242 9154 14254
rect 16046 14306 16098 14318
rect 16046 14242 16098 14254
rect 17950 14306 18002 14318
rect 17950 14242 18002 14254
rect 18510 14306 18562 14318
rect 18510 14242 18562 14254
rect 23998 14306 24050 14318
rect 23998 14242 24050 14254
rect 24222 14306 24274 14318
rect 24222 14242 24274 14254
rect 26126 14306 26178 14318
rect 26126 14242 26178 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 31502 14306 31554 14318
rect 46846 14306 46898 14318
rect 46498 14254 46510 14306
rect 46562 14254 46574 14306
rect 31502 14242 31554 14254
rect 46846 14242 46898 14254
rect 47406 14306 47458 14318
rect 47406 14242 47458 14254
rect 51438 14306 51490 14318
rect 51438 14242 51490 14254
rect 53230 14306 53282 14318
rect 53230 14242 53282 14254
rect 1344 14138 53648 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 53648 14138
rect 1344 14052 53648 14086
rect 5854 13970 5906 13982
rect 5854 13906 5906 13918
rect 7310 13970 7362 13982
rect 7310 13906 7362 13918
rect 7422 13970 7474 13982
rect 7422 13906 7474 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 10110 13970 10162 13982
rect 10110 13906 10162 13918
rect 12686 13970 12738 13982
rect 12686 13906 12738 13918
rect 13134 13970 13186 13982
rect 13134 13906 13186 13918
rect 40014 13970 40066 13982
rect 40014 13906 40066 13918
rect 46398 13970 46450 13982
rect 46398 13906 46450 13918
rect 53342 13970 53394 13982
rect 53342 13906 53394 13918
rect 7534 13858 7586 13870
rect 5282 13806 5294 13858
rect 5346 13806 5358 13858
rect 7534 13794 7586 13806
rect 8766 13858 8818 13870
rect 8766 13794 8818 13806
rect 8878 13858 8930 13870
rect 10894 13858 10946 13870
rect 10434 13806 10446 13858
rect 10498 13806 10510 13858
rect 8878 13794 8930 13806
rect 10894 13794 10946 13806
rect 11230 13858 11282 13870
rect 11230 13794 11282 13806
rect 11566 13858 11618 13870
rect 20974 13858 21026 13870
rect 40126 13858 40178 13870
rect 12338 13806 12350 13858
rect 12402 13806 12414 13858
rect 39330 13806 39342 13858
rect 39394 13806 39406 13858
rect 46722 13806 46734 13858
rect 46786 13806 46798 13858
rect 11566 13794 11618 13806
rect 20974 13794 21026 13806
rect 40126 13794 40178 13806
rect 4958 13746 5010 13758
rect 7982 13746 8034 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 5618 13694 5630 13746
rect 5682 13694 5694 13746
rect 4958 13682 5010 13694
rect 7982 13682 8034 13694
rect 8654 13746 8706 13758
rect 25790 13746 25842 13758
rect 11890 13694 11902 13746
rect 11954 13694 11966 13746
rect 24658 13694 24670 13746
rect 24722 13694 24734 13746
rect 8654 13682 8706 13694
rect 25790 13682 25842 13694
rect 26014 13746 26066 13758
rect 26014 13682 26066 13694
rect 26350 13746 26402 13758
rect 36654 13746 36706 13758
rect 26562 13694 26574 13746
rect 26626 13694 26638 13746
rect 36082 13694 36094 13746
rect 36146 13694 36158 13746
rect 26350 13682 26402 13694
rect 36654 13682 36706 13694
rect 38558 13746 38610 13758
rect 39902 13746 39954 13758
rect 39106 13694 39118 13746
rect 39170 13694 39182 13746
rect 39666 13694 39678 13746
rect 39730 13694 39742 13746
rect 38558 13682 38610 13694
rect 39902 13682 39954 13694
rect 40238 13746 40290 13758
rect 45166 13746 45218 13758
rect 44706 13694 44718 13746
rect 44770 13694 44782 13746
rect 40238 13682 40290 13694
rect 45166 13682 45218 13694
rect 25342 13634 25394 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 11778 13582 11790 13634
rect 11842 13582 11854 13634
rect 21746 13582 21758 13634
rect 21810 13582 21822 13634
rect 23874 13582 23886 13634
rect 23938 13582 23950 13634
rect 25342 13570 25394 13582
rect 26126 13634 26178 13646
rect 27346 13582 27358 13634
rect 27410 13582 27422 13634
rect 29474 13582 29486 13634
rect 29538 13582 29550 13634
rect 35746 13582 35758 13634
rect 35810 13582 35822 13634
rect 41794 13582 41806 13634
rect 41858 13582 41870 13634
rect 43922 13582 43934 13634
rect 43986 13582 43998 13634
rect 26126 13570 26178 13582
rect 5966 13522 6018 13534
rect 20862 13522 20914 13534
rect 8194 13470 8206 13522
rect 8258 13470 8270 13522
rect 5966 13458 6018 13470
rect 20862 13458 20914 13470
rect 38670 13522 38722 13534
rect 38670 13458 38722 13470
rect 1344 13354 53648 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 53648 13354
rect 1344 13268 53648 13302
rect 15934 13186 15986 13198
rect 15934 13122 15986 13134
rect 17614 13186 17666 13198
rect 17614 13122 17666 13134
rect 18286 13186 18338 13198
rect 18286 13122 18338 13134
rect 37886 13186 37938 13198
rect 37886 13122 37938 13134
rect 42590 13186 42642 13198
rect 42590 13122 42642 13134
rect 10782 13074 10834 13086
rect 10782 13010 10834 13022
rect 12238 13074 12290 13086
rect 12238 13010 12290 13022
rect 14590 13074 14642 13086
rect 14590 13010 14642 13022
rect 19070 13074 19122 13086
rect 35422 13074 35474 13086
rect 24098 13022 24110 13074
rect 24162 13022 24174 13074
rect 33618 13022 33630 13074
rect 33682 13022 33694 13074
rect 19070 13010 19122 13022
rect 35422 13010 35474 13022
rect 37550 13074 37602 13086
rect 43038 13074 43090 13086
rect 41010 13022 41022 13074
rect 41074 13022 41086 13074
rect 37550 13010 37602 13022
rect 43038 13010 43090 13022
rect 2606 12962 2658 12974
rect 2606 12898 2658 12910
rect 8542 12962 8594 12974
rect 16382 12962 16434 12974
rect 11442 12910 11454 12962
rect 11506 12910 11518 12962
rect 15586 12910 15598 12962
rect 15650 12910 15662 12962
rect 8542 12898 8594 12910
rect 16382 12898 16434 12910
rect 17166 12962 17218 12974
rect 18398 12962 18450 12974
rect 26350 12962 26402 12974
rect 17378 12910 17390 12962
rect 17442 12910 17454 12962
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 26114 12910 26126 12962
rect 26178 12910 26190 12962
rect 17166 12898 17218 12910
rect 18398 12898 18450 12910
rect 26350 12898 26402 12910
rect 26686 12962 26738 12974
rect 38670 12962 38722 12974
rect 40910 12962 40962 12974
rect 30706 12910 30718 12962
rect 30770 12910 30782 12962
rect 35970 12910 35982 12962
rect 36034 12910 36046 12962
rect 38210 12910 38222 12962
rect 38274 12910 38286 12962
rect 39106 12910 39118 12962
rect 39170 12910 39182 12962
rect 26686 12898 26738 12910
rect 38670 12898 38722 12910
rect 40910 12898 40962 12910
rect 42254 12962 42306 12974
rect 42254 12898 42306 12910
rect 2270 12850 2322 12862
rect 2270 12786 2322 12798
rect 8430 12850 8482 12862
rect 16830 12850 16882 12862
rect 34638 12850 34690 12862
rect 35758 12850 35810 12862
rect 13794 12798 13806 12850
rect 13858 12798 13870 12850
rect 16146 12798 16158 12850
rect 16210 12798 16222 12850
rect 31490 12798 31502 12850
rect 31554 12798 31566 12850
rect 35522 12798 35534 12850
rect 35586 12798 35598 12850
rect 8430 12786 8482 12798
rect 16830 12786 16882 12798
rect 34638 12786 34690 12798
rect 35758 12786 35810 12798
rect 39566 12850 39618 12862
rect 39566 12786 39618 12798
rect 40462 12850 40514 12862
rect 40462 12786 40514 12798
rect 42478 12850 42530 12862
rect 42478 12786 42530 12798
rect 4846 12738 4898 12750
rect 4846 12674 4898 12686
rect 8206 12738 8258 12750
rect 8206 12674 8258 12686
rect 11230 12738 11282 12750
rect 11230 12674 11282 12686
rect 13470 12738 13522 12750
rect 26574 12738 26626 12750
rect 15922 12686 15934 12738
rect 15986 12686 15998 12738
rect 17602 12686 17614 12738
rect 17666 12686 17678 12738
rect 13470 12674 13522 12686
rect 26574 12674 26626 12686
rect 27134 12738 27186 12750
rect 36430 12738 36482 12750
rect 34290 12686 34302 12738
rect 34354 12686 34366 12738
rect 27134 12674 27186 12686
rect 36430 12674 36482 12686
rect 37998 12738 38050 12750
rect 37998 12674 38050 12686
rect 40686 12738 40738 12750
rect 40686 12674 40738 12686
rect 41022 12738 41074 12750
rect 41022 12674 41074 12686
rect 1344 12570 53648 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 53648 12570
rect 1344 12484 53648 12518
rect 7758 12402 7810 12414
rect 7758 12338 7810 12350
rect 7870 12402 7922 12414
rect 7870 12338 7922 12350
rect 8430 12402 8482 12414
rect 8430 12338 8482 12350
rect 15150 12402 15202 12414
rect 15150 12338 15202 12350
rect 19966 12402 20018 12414
rect 19966 12338 20018 12350
rect 23886 12402 23938 12414
rect 23886 12338 23938 12350
rect 28254 12402 28306 12414
rect 28254 12338 28306 12350
rect 31838 12402 31890 12414
rect 31838 12338 31890 12350
rect 35086 12402 35138 12414
rect 35086 12338 35138 12350
rect 35310 12402 35362 12414
rect 35310 12338 35362 12350
rect 35422 12402 35474 12414
rect 35422 12338 35474 12350
rect 36094 12402 36146 12414
rect 36094 12338 36146 12350
rect 36206 12402 36258 12414
rect 36206 12338 36258 12350
rect 38670 12402 38722 12414
rect 38670 12338 38722 12350
rect 44606 12402 44658 12414
rect 44606 12338 44658 12350
rect 44942 12402 44994 12414
rect 44942 12338 44994 12350
rect 46062 12402 46114 12414
rect 46062 12338 46114 12350
rect 49870 12402 49922 12414
rect 49870 12338 49922 12350
rect 5966 12290 6018 12302
rect 14366 12290 14418 12302
rect 7074 12238 7086 12290
rect 7138 12238 7150 12290
rect 14130 12238 14142 12290
rect 14194 12238 14206 12290
rect 5966 12226 6018 12238
rect 14366 12226 14418 12238
rect 14926 12290 14978 12302
rect 14926 12226 14978 12238
rect 17390 12290 17442 12302
rect 17390 12226 17442 12238
rect 23550 12290 23602 12302
rect 23550 12226 23602 12238
rect 24110 12290 24162 12302
rect 24110 12226 24162 12238
rect 24558 12290 24610 12302
rect 24558 12226 24610 12238
rect 36318 12290 36370 12302
rect 38994 12238 39006 12290
rect 39058 12238 39070 12290
rect 51090 12238 51102 12290
rect 51154 12238 51166 12290
rect 36318 12226 36370 12238
rect 6414 12178 6466 12190
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 6414 12114 6466 12126
rect 6638 12178 6690 12190
rect 6638 12114 6690 12126
rect 6862 12178 6914 12190
rect 6862 12114 6914 12126
rect 7422 12178 7474 12190
rect 13918 12178 13970 12190
rect 13570 12126 13582 12178
rect 13634 12126 13646 12178
rect 7422 12114 7474 12126
rect 13918 12114 13970 12126
rect 15598 12178 15650 12190
rect 16046 12178 16098 12190
rect 17838 12178 17890 12190
rect 23774 12178 23826 12190
rect 15810 12126 15822 12178
rect 15874 12126 15886 12178
rect 16370 12126 16382 12178
rect 16434 12126 16446 12178
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 18050 12126 18062 12178
rect 18114 12126 18126 12178
rect 15598 12114 15650 12126
rect 16046 12114 16098 12126
rect 17838 12114 17890 12126
rect 23774 12114 23826 12126
rect 24334 12178 24386 12190
rect 24334 12114 24386 12126
rect 24670 12178 24722 12190
rect 34750 12178 34802 12190
rect 25778 12126 25790 12178
rect 25842 12126 25854 12178
rect 32050 12126 32062 12178
rect 32114 12126 32126 12178
rect 24670 12114 24722 12126
rect 34750 12114 34802 12126
rect 35870 12178 35922 12190
rect 35870 12114 35922 12126
rect 35982 12178 36034 12190
rect 35982 12114 36034 12126
rect 38110 12178 38162 12190
rect 38110 12114 38162 12126
rect 38334 12178 38386 12190
rect 38334 12114 38386 12126
rect 44830 12178 44882 12190
rect 44830 12114 44882 12126
rect 45054 12178 45106 12190
rect 45054 12114 45106 12126
rect 49534 12178 49586 12190
rect 50306 12126 50318 12178
rect 50370 12126 50382 12178
rect 49534 12114 49586 12126
rect 6078 12066 6130 12078
rect 5394 12014 5406 12066
rect 5458 12014 5470 12066
rect 6078 12002 6130 12014
rect 6526 12066 6578 12078
rect 6526 12002 6578 12014
rect 14254 12066 14306 12078
rect 15710 12066 15762 12078
rect 15250 12014 15262 12066
rect 15314 12014 15326 12066
rect 14254 12002 14306 12014
rect 15710 12002 15762 12014
rect 17502 12066 17554 12078
rect 49198 12066 49250 12078
rect 20402 12014 20414 12066
rect 20466 12014 20478 12066
rect 26898 12014 26910 12066
rect 26962 12014 26974 12066
rect 53218 12014 53230 12066
rect 53282 12014 53294 12066
rect 17502 12002 17554 12014
rect 49198 12002 49250 12014
rect 5182 11954 5234 11966
rect 5182 11890 5234 11902
rect 7646 11954 7698 11966
rect 7646 11890 7698 11902
rect 31726 11954 31778 11966
rect 37762 11902 37774 11954
rect 37826 11902 37838 11954
rect 31726 11890 31778 11902
rect 1344 11786 53648 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 53648 11786
rect 1344 11700 53648 11734
rect 6190 11618 6242 11630
rect 6190 11554 6242 11566
rect 9102 11618 9154 11630
rect 9102 11554 9154 11566
rect 9326 11618 9378 11630
rect 9326 11554 9378 11566
rect 11118 11618 11170 11630
rect 23214 11618 23266 11630
rect 13682 11566 13694 11618
rect 13746 11566 13758 11618
rect 11118 11554 11170 11566
rect 23214 11554 23266 11566
rect 6414 11506 6466 11518
rect 17726 11506 17778 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 15810 11454 15822 11506
rect 15874 11454 15886 11506
rect 6414 11442 6466 11454
rect 17726 11442 17778 11454
rect 21422 11506 21474 11518
rect 21422 11442 21474 11454
rect 27918 11506 27970 11518
rect 27918 11442 27970 11454
rect 31726 11506 31778 11518
rect 31726 11442 31778 11454
rect 32510 11506 32562 11518
rect 49074 11454 49086 11506
rect 49138 11454 49150 11506
rect 32510 11442 32562 11454
rect 5742 11394 5794 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 5742 11330 5794 11342
rect 8878 11394 8930 11406
rect 12798 11394 12850 11406
rect 26574 11394 26626 11406
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 14018 11342 14030 11394
rect 14082 11342 14094 11394
rect 15250 11342 15262 11394
rect 15314 11342 15326 11394
rect 20402 11342 20414 11394
rect 20466 11342 20478 11394
rect 8878 11330 8930 11342
rect 12798 11330 12850 11342
rect 26574 11330 26626 11342
rect 27022 11394 27074 11406
rect 29262 11394 29314 11406
rect 30942 11394 30994 11406
rect 27346 11342 27358 11394
rect 27410 11342 27422 11394
rect 29474 11342 29486 11394
rect 29538 11342 29550 11394
rect 27022 11330 27074 11342
rect 29262 11330 29314 11342
rect 30942 11330 30994 11342
rect 31166 11394 31218 11406
rect 31166 11330 31218 11342
rect 31614 11394 31666 11406
rect 32622 11394 32674 11406
rect 45166 11394 45218 11406
rect 32162 11342 32174 11394
rect 32226 11342 32238 11394
rect 32834 11342 32846 11394
rect 32898 11342 32910 11394
rect 40786 11342 40798 11394
rect 40850 11342 40862 11394
rect 41458 11342 41470 11394
rect 41522 11342 41534 11394
rect 31614 11330 31666 11342
rect 32622 11330 32674 11342
rect 45166 11330 45218 11342
rect 45838 11394 45890 11406
rect 46274 11342 46286 11394
rect 46338 11342 46350 11394
rect 46946 11342 46958 11394
rect 47010 11342 47022 11394
rect 45838 11330 45890 11342
rect 5630 11282 5682 11294
rect 5630 11218 5682 11230
rect 10670 11282 10722 11294
rect 12910 11282 12962 11294
rect 10882 11230 10894 11282
rect 10946 11230 10958 11282
rect 10670 11218 10722 11230
rect 12910 11218 12962 11230
rect 14254 11282 14306 11294
rect 14254 11218 14306 11230
rect 20750 11282 20802 11294
rect 20750 11218 20802 11230
rect 23326 11282 23378 11294
rect 29150 11282 29202 11294
rect 25890 11230 25902 11282
rect 25954 11230 25966 11282
rect 26786 11230 26798 11282
rect 26850 11230 26862 11282
rect 23326 11218 23378 11230
rect 29150 11218 29202 11230
rect 45950 11282 46002 11294
rect 45950 11218 46002 11230
rect 50654 11282 50706 11294
rect 50654 11218 50706 11230
rect 52222 11282 52274 11294
rect 52222 11218 52274 11230
rect 52894 11282 52946 11294
rect 52894 11218 52946 11230
rect 53230 11282 53282 11294
rect 53230 11218 53282 11230
rect 5070 11170 5122 11182
rect 5070 11106 5122 11118
rect 6526 11170 6578 11182
rect 6526 11106 6578 11118
rect 9774 11170 9826 11182
rect 12686 11170 12738 11182
rect 11106 11118 11118 11170
rect 11170 11118 11182 11170
rect 9774 11106 9826 11118
rect 12686 11106 12738 11118
rect 13470 11170 13522 11182
rect 13470 11106 13522 11118
rect 20638 11170 20690 11182
rect 20638 11106 20690 11118
rect 23214 11170 23266 11182
rect 23214 11106 23266 11118
rect 24334 11170 24386 11182
rect 24334 11106 24386 11118
rect 26238 11170 26290 11182
rect 26238 11106 26290 11118
rect 27358 11170 27410 11182
rect 27358 11106 27410 11118
rect 31838 11170 31890 11182
rect 31838 11106 31890 11118
rect 32398 11170 32450 11182
rect 42366 11170 42418 11182
rect 41010 11118 41022 11170
rect 41074 11118 41086 11170
rect 41682 11118 41694 11170
rect 41746 11118 41758 11170
rect 42018 11118 42030 11170
rect 42082 11118 42094 11170
rect 32398 11106 32450 11118
rect 42366 11106 42418 11118
rect 42814 11170 42866 11182
rect 42814 11106 42866 11118
rect 43262 11170 43314 11182
rect 43262 11106 43314 11118
rect 45390 11170 45442 11182
rect 45390 11106 45442 11118
rect 45614 11170 45666 11182
rect 45614 11106 45666 11118
rect 49534 11170 49586 11182
rect 49534 11106 49586 11118
rect 49982 11170 50034 11182
rect 49982 11106 50034 11118
rect 50766 11170 50818 11182
rect 50766 11106 50818 11118
rect 1344 11002 53648 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 53648 11002
rect 1344 10916 53648 10950
rect 10334 10834 10386 10846
rect 10334 10770 10386 10782
rect 17502 10834 17554 10846
rect 17502 10770 17554 10782
rect 18734 10834 18786 10846
rect 18734 10770 18786 10782
rect 19630 10834 19682 10846
rect 19630 10770 19682 10782
rect 23774 10834 23826 10846
rect 23774 10770 23826 10782
rect 23886 10834 23938 10846
rect 30942 10834 30994 10846
rect 30370 10782 30382 10834
rect 30434 10782 30446 10834
rect 23886 10770 23938 10782
rect 30942 10770 30994 10782
rect 31950 10834 32002 10846
rect 31950 10770 32002 10782
rect 32174 10834 32226 10846
rect 32174 10770 32226 10782
rect 37326 10834 37378 10846
rect 37326 10770 37378 10782
rect 40462 10834 40514 10846
rect 40462 10770 40514 10782
rect 41358 10834 41410 10846
rect 41358 10770 41410 10782
rect 41918 10834 41970 10846
rect 45602 10782 45614 10834
rect 45666 10782 45678 10834
rect 49634 10782 49646 10834
rect 49698 10782 49710 10834
rect 41918 10770 41970 10782
rect 9550 10722 9602 10734
rect 9550 10658 9602 10670
rect 9886 10722 9938 10734
rect 9886 10658 9938 10670
rect 10558 10722 10610 10734
rect 13694 10722 13746 10734
rect 11442 10670 11454 10722
rect 11506 10670 11518 10722
rect 10558 10658 10610 10670
rect 13694 10658 13746 10670
rect 13918 10722 13970 10734
rect 23438 10722 23490 10734
rect 20738 10670 20750 10722
rect 20802 10670 20814 10722
rect 13918 10658 13970 10670
rect 23438 10658 23490 10670
rect 23550 10722 23602 10734
rect 23550 10658 23602 10670
rect 24110 10722 24162 10734
rect 24110 10658 24162 10670
rect 24222 10722 24274 10734
rect 31838 10722 31890 10734
rect 36766 10722 36818 10734
rect 39454 10722 39506 10734
rect 25218 10670 25230 10722
rect 25282 10670 25294 10722
rect 27570 10670 27582 10722
rect 27634 10670 27646 10722
rect 36418 10670 36430 10722
rect 36482 10670 36494 10722
rect 38994 10670 39006 10722
rect 39058 10670 39070 10722
rect 24222 10658 24274 10670
rect 31838 10658 31890 10670
rect 36766 10658 36818 10670
rect 39454 10658 39506 10670
rect 39566 10722 39618 10734
rect 39566 10658 39618 10670
rect 42142 10722 42194 10734
rect 51090 10670 51102 10722
rect 51154 10670 51166 10722
rect 42142 10658 42194 10670
rect 5742 10610 5794 10622
rect 5742 10546 5794 10558
rect 6078 10610 6130 10622
rect 6078 10546 6130 10558
rect 6302 10610 6354 10622
rect 6302 10546 6354 10558
rect 6638 10610 6690 10622
rect 6638 10546 6690 10558
rect 7086 10610 7138 10622
rect 7086 10546 7138 10558
rect 10110 10610 10162 10622
rect 10110 10546 10162 10558
rect 10670 10610 10722 10622
rect 10670 10546 10722 10558
rect 11118 10610 11170 10622
rect 25566 10610 25618 10622
rect 35646 10610 35698 10622
rect 16818 10558 16830 10610
rect 16882 10558 16894 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 26898 10558 26910 10610
rect 26962 10558 26974 10610
rect 30146 10558 30158 10610
rect 30210 10558 30222 10610
rect 11118 10546 11170 10558
rect 25566 10546 25618 10558
rect 35646 10546 35698 10558
rect 35870 10610 35922 10622
rect 35870 10546 35922 10558
rect 36206 10610 36258 10622
rect 41134 10610 41186 10622
rect 38770 10558 38782 10610
rect 38834 10558 38846 10610
rect 36206 10546 36258 10558
rect 41134 10546 41186 10558
rect 41470 10610 41522 10622
rect 43822 10610 43874 10622
rect 42914 10558 42926 10610
rect 42978 10558 42990 10610
rect 43362 10558 43374 10610
rect 43426 10558 43438 10610
rect 41470 10546 41522 10558
rect 43822 10546 43874 10558
rect 45166 10610 45218 10622
rect 49198 10610 49250 10622
rect 49646 10610 49698 10622
rect 45378 10558 45390 10610
rect 45442 10558 45454 10610
rect 49410 10558 49422 10610
rect 49474 10558 49486 10610
rect 49858 10558 49870 10610
rect 49922 10558 49934 10610
rect 50306 10558 50318 10610
rect 50370 10558 50382 10610
rect 45166 10546 45218 10558
rect 49198 10546 49250 10558
rect 49646 10546 49698 10558
rect 5630 10498 5682 10510
rect 5630 10434 5682 10446
rect 6190 10498 6242 10510
rect 6190 10434 6242 10446
rect 7422 10498 7474 10510
rect 7422 10434 7474 10446
rect 9662 10498 9714 10510
rect 18846 10498 18898 10510
rect 26014 10498 26066 10510
rect 35982 10498 36034 10510
rect 13570 10446 13582 10498
rect 13634 10446 13646 10498
rect 15698 10446 15710 10498
rect 15762 10446 15774 10498
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 29698 10446 29710 10498
rect 29762 10446 29774 10498
rect 41906 10446 41918 10498
rect 41970 10446 41982 10498
rect 45042 10446 45054 10498
rect 45106 10446 45118 10498
rect 53218 10446 53230 10498
rect 53282 10446 53294 10498
rect 9662 10434 9714 10446
rect 18846 10434 18898 10446
rect 26014 10434 26066 10446
rect 35982 10434 36034 10446
rect 6526 10386 6578 10398
rect 6526 10322 6578 10334
rect 39678 10386 39730 10398
rect 43922 10334 43934 10386
rect 43986 10334 43998 10386
rect 39678 10322 39730 10334
rect 1344 10218 53648 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 53648 10218
rect 1344 10132 53648 10166
rect 12462 10050 12514 10062
rect 11218 9998 11230 10050
rect 11282 9998 11294 10050
rect 12462 9986 12514 9998
rect 14030 10050 14082 10062
rect 14030 9986 14082 9998
rect 23550 10050 23602 10062
rect 23550 9986 23602 9998
rect 27246 10050 27298 10062
rect 27246 9986 27298 9998
rect 39230 10050 39282 10062
rect 39230 9986 39282 9998
rect 44942 10050 44994 10062
rect 44942 9986 44994 9998
rect 47406 10050 47458 10062
rect 47406 9986 47458 9998
rect 10446 9938 10498 9950
rect 2146 9886 2158 9938
rect 2210 9886 2222 9938
rect 4274 9886 4286 9938
rect 4338 9886 4350 9938
rect 10446 9874 10498 9886
rect 15038 9938 15090 9950
rect 29934 9938 29986 9950
rect 17378 9886 17390 9938
rect 17442 9886 17454 9938
rect 19506 9886 19518 9938
rect 19570 9886 19582 9938
rect 15038 9874 15090 9886
rect 29934 9874 29986 9886
rect 11790 9826 11842 9838
rect 12910 9826 12962 9838
rect 14478 9826 14530 9838
rect 23662 9826 23714 9838
rect 5058 9774 5070 9826
rect 5122 9774 5134 9826
rect 11106 9774 11118 9826
rect 11170 9774 11182 9826
rect 11554 9774 11566 9826
rect 11618 9774 11630 9826
rect 12338 9774 12350 9826
rect 12402 9774 12414 9826
rect 13906 9774 13918 9826
rect 13970 9774 13982 9826
rect 16594 9774 16606 9826
rect 16658 9774 16670 9826
rect 11790 9762 11842 9774
rect 12910 9762 12962 9774
rect 14478 9762 14530 9774
rect 23662 9762 23714 9774
rect 27134 9826 27186 9838
rect 27134 9762 27186 9774
rect 29486 9826 29538 9838
rect 36206 9826 36258 9838
rect 33842 9774 33854 9826
rect 33906 9774 33918 9826
rect 29486 9762 29538 9774
rect 36206 9762 36258 9774
rect 38446 9826 38498 9838
rect 38446 9762 38498 9774
rect 38670 9826 38722 9838
rect 38670 9762 38722 9774
rect 39118 9826 39170 9838
rect 45390 9826 45442 9838
rect 41346 9774 41358 9826
rect 41410 9774 41422 9826
rect 41794 9774 41806 9826
rect 41858 9774 41870 9826
rect 39118 9762 39170 9774
rect 45390 9762 45442 9774
rect 45614 9826 45666 9838
rect 45614 9762 45666 9774
rect 45838 9826 45890 9838
rect 45838 9762 45890 9774
rect 46398 9826 46450 9838
rect 46398 9762 46450 9774
rect 46846 9826 46898 9838
rect 48414 9826 48466 9838
rect 47842 9774 47854 9826
rect 47906 9774 47918 9826
rect 46846 9762 46898 9774
rect 48414 9762 48466 9774
rect 36094 9714 36146 9726
rect 12674 9662 12686 9714
rect 12738 9662 12750 9714
rect 14242 9662 14254 9714
rect 14306 9662 14318 9714
rect 29138 9662 29150 9714
rect 29202 9662 29214 9714
rect 36094 9650 36146 9662
rect 38894 9714 38946 9726
rect 38894 9650 38946 9662
rect 40910 9714 40962 9726
rect 46062 9714 46114 9726
rect 43586 9662 43598 9714
rect 43650 9662 43662 9714
rect 40910 9650 40962 9662
rect 46062 9650 46114 9662
rect 48078 9714 48130 9726
rect 48078 9650 48130 9662
rect 48190 9714 48242 9726
rect 49870 9714 49922 9726
rect 50542 9714 50594 9726
rect 49522 9662 49534 9714
rect 49586 9662 49598 9714
rect 50194 9662 50206 9714
rect 50258 9662 50270 9714
rect 48190 9650 48242 9662
rect 49870 9650 49922 9662
rect 50542 9650 50594 9662
rect 5742 9602 5794 9614
rect 5742 9538 5794 9550
rect 11006 9602 11058 9614
rect 11006 9538 11058 9550
rect 12126 9602 12178 9614
rect 15374 9602 15426 9614
rect 14130 9550 14142 9602
rect 14194 9550 14206 9602
rect 12126 9538 12178 9550
rect 15374 9538 15426 9550
rect 16270 9602 16322 9614
rect 16270 9538 16322 9550
rect 23550 9602 23602 9614
rect 23550 9538 23602 9550
rect 27246 9602 27298 9614
rect 35870 9602 35922 9614
rect 46510 9602 46562 9614
rect 33618 9550 33630 9602
rect 33682 9550 33694 9602
rect 40786 9550 40798 9602
rect 40850 9550 40862 9602
rect 27246 9538 27298 9550
rect 35870 9538 35922 9550
rect 46510 9538 46562 9550
rect 1344 9434 53648 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 53648 9434
rect 1344 9348 53648 9382
rect 12126 9266 12178 9278
rect 12126 9202 12178 9214
rect 13246 9266 13298 9278
rect 13246 9202 13298 9214
rect 16718 9266 16770 9278
rect 16718 9202 16770 9214
rect 26238 9266 26290 9278
rect 26238 9202 26290 9214
rect 29822 9266 29874 9278
rect 35646 9266 35698 9278
rect 31714 9214 31726 9266
rect 31778 9214 31790 9266
rect 29822 9202 29874 9214
rect 35646 9202 35698 9214
rect 36430 9266 36482 9278
rect 36430 9202 36482 9214
rect 38334 9266 38386 9278
rect 38334 9202 38386 9214
rect 42254 9266 42306 9278
rect 42254 9202 42306 9214
rect 43822 9266 43874 9278
rect 43822 9202 43874 9214
rect 23438 9154 23490 9166
rect 32174 9154 32226 9166
rect 23762 9102 23774 9154
rect 23826 9102 23838 9154
rect 31938 9102 31950 9154
rect 32002 9102 32014 9154
rect 23438 9090 23490 9102
rect 32174 9090 32226 9102
rect 33406 9154 33458 9166
rect 33406 9090 33458 9102
rect 35870 9154 35922 9166
rect 35870 9090 35922 9102
rect 36878 9154 36930 9166
rect 36878 9090 36930 9102
rect 38110 9154 38162 9166
rect 38110 9090 38162 9102
rect 29262 9042 29314 9054
rect 29262 8978 29314 8990
rect 31054 9042 31106 9054
rect 35422 9042 35474 9054
rect 31378 8990 31390 9042
rect 31442 8990 31454 9042
rect 33058 8990 33070 9042
rect 33122 8990 33134 9042
rect 35186 8990 35198 9042
rect 35250 8990 35262 9042
rect 31054 8978 31106 8990
rect 35422 8978 35474 8990
rect 36318 9042 36370 9054
rect 36318 8978 36370 8990
rect 36654 9042 36706 9054
rect 36654 8978 36706 8990
rect 42142 9042 42194 9054
rect 42142 8978 42194 8990
rect 42478 9042 42530 9054
rect 42478 8978 42530 8990
rect 45166 9042 45218 9054
rect 45166 8978 45218 8990
rect 45390 9042 45442 9054
rect 45390 8978 45442 8990
rect 45838 9042 45890 9054
rect 52782 9042 52834 9054
rect 52210 8990 52222 9042
rect 52274 8990 52286 9042
rect 45838 8978 45890 8990
rect 52782 8978 52834 8990
rect 16830 8930 16882 8942
rect 16830 8866 16882 8878
rect 26126 8930 26178 8942
rect 42814 8930 42866 8942
rect 35298 8878 35310 8930
rect 35362 8878 35374 8930
rect 38434 8878 38446 8930
rect 38498 8878 38510 8930
rect 45714 8878 45726 8930
rect 45778 8878 45790 8930
rect 26126 8866 26178 8878
rect 42814 8866 42866 8878
rect 31726 8818 31778 8830
rect 31726 8754 31778 8766
rect 33070 8818 33122 8830
rect 33070 8754 33122 8766
rect 36766 8818 36818 8830
rect 36766 8754 36818 8766
rect 45950 8818 46002 8830
rect 45950 8754 46002 8766
rect 52558 8818 52610 8830
rect 52558 8754 52610 8766
rect 1344 8650 53648 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 53648 8650
rect 1344 8564 53648 8598
rect 12798 8482 12850 8494
rect 12798 8418 12850 8430
rect 47294 8482 47346 8494
rect 47294 8418 47346 8430
rect 26238 8370 26290 8382
rect 8082 8318 8094 8370
rect 8146 8318 8158 8370
rect 10210 8318 10222 8370
rect 10274 8318 10286 8370
rect 15362 8318 15374 8370
rect 15426 8318 15438 8370
rect 17490 8318 17502 8370
rect 17554 8318 17566 8370
rect 22978 8318 22990 8370
rect 23042 8318 23054 8370
rect 25330 8318 25342 8370
rect 25394 8318 25406 8370
rect 26238 8306 26290 8318
rect 27246 8370 27298 8382
rect 36318 8370 36370 8382
rect 31602 8318 31614 8370
rect 31666 8318 31678 8370
rect 33730 8318 33742 8370
rect 33794 8318 33806 8370
rect 39330 8318 39342 8370
rect 39394 8318 39406 8370
rect 27246 8306 27298 8318
rect 36318 8306 36370 8318
rect 20638 8258 20690 8270
rect 7410 8206 7422 8258
rect 7474 8206 7486 8258
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 19730 8206 19742 8258
rect 19794 8206 19806 8258
rect 20290 8206 20302 8258
rect 20354 8206 20366 8258
rect 20638 8194 20690 8206
rect 25230 8258 25282 8270
rect 26014 8258 26066 8270
rect 35646 8258 35698 8270
rect 25442 8206 25454 8258
rect 25506 8206 25518 8258
rect 26674 8206 26686 8258
rect 26738 8206 26750 8258
rect 30818 8206 30830 8258
rect 30882 8206 30894 8258
rect 25230 8194 25282 8206
rect 26014 8194 26066 8206
rect 35646 8194 35698 8206
rect 35870 8258 35922 8270
rect 38894 8258 38946 8270
rect 37202 8206 37214 8258
rect 37266 8206 37278 8258
rect 35870 8194 35922 8206
rect 38894 8194 38946 8206
rect 41470 8258 41522 8270
rect 41470 8194 41522 8206
rect 42702 8258 42754 8270
rect 42702 8194 42754 8206
rect 42926 8258 42978 8270
rect 42926 8194 42978 8206
rect 43150 8258 43202 8270
rect 53230 8258 53282 8270
rect 43922 8206 43934 8258
rect 43986 8206 43998 8258
rect 47170 8206 47182 8258
rect 47234 8206 47246 8258
rect 49074 8206 49086 8258
rect 49138 8206 49150 8258
rect 43150 8194 43202 8206
rect 53230 8194 53282 8206
rect 12910 8146 12962 8158
rect 12910 8082 12962 8094
rect 23550 8146 23602 8158
rect 23550 8082 23602 8094
rect 24782 8146 24834 8158
rect 24782 8082 24834 8094
rect 25790 8146 25842 8158
rect 34750 8146 34802 8158
rect 26450 8094 26462 8146
rect 26514 8094 26526 8146
rect 25790 8082 25842 8094
rect 34750 8082 34802 8094
rect 34974 8146 35026 8158
rect 34974 8082 35026 8094
rect 35422 8146 35474 8158
rect 35422 8082 35474 8094
rect 35758 8146 35810 8158
rect 39454 8146 39506 8158
rect 36978 8094 36990 8146
rect 37042 8094 37054 8146
rect 35758 8082 35810 8094
rect 39454 8082 39506 8094
rect 41806 8146 41858 8158
rect 41806 8082 41858 8094
rect 43374 8146 43426 8158
rect 48626 8094 48638 8146
rect 48690 8094 48702 8146
rect 49746 8094 49758 8146
rect 49810 8094 49822 8146
rect 52882 8094 52894 8146
rect 52946 8094 52958 8146
rect 43374 8082 43426 8094
rect 10670 8034 10722 8046
rect 10670 7970 10722 7982
rect 17950 8034 18002 8046
rect 20526 8034 20578 8046
rect 19506 7982 19518 8034
rect 19570 7982 19582 8034
rect 17950 7970 18002 7982
rect 20526 7970 20578 7982
rect 22990 8034 23042 8046
rect 22990 7970 23042 7982
rect 23102 8034 23154 8046
rect 23102 7970 23154 7982
rect 23326 8034 23378 8046
rect 23326 7970 23378 7982
rect 25006 8034 25058 8046
rect 34862 8034 34914 8046
rect 26338 7982 26350 8034
rect 26402 7982 26414 8034
rect 25006 7970 25058 7982
rect 34862 7970 34914 7982
rect 39230 8034 39282 8046
rect 39230 7970 39282 7982
rect 42590 8034 42642 8046
rect 43698 7982 43710 8034
rect 43762 7982 43774 8034
rect 42590 7970 42642 7982
rect 1344 7866 53648 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 53648 7866
rect 1344 7780 53648 7814
rect 23102 7698 23154 7710
rect 23102 7634 23154 7646
rect 23326 7698 23378 7710
rect 23326 7634 23378 7646
rect 25902 7698 25954 7710
rect 25902 7634 25954 7646
rect 31166 7698 31218 7710
rect 31166 7634 31218 7646
rect 31838 7698 31890 7710
rect 31838 7634 31890 7646
rect 39006 7698 39058 7710
rect 39006 7634 39058 7646
rect 40910 7698 40962 7710
rect 40910 7634 40962 7646
rect 42142 7698 42194 7710
rect 42142 7634 42194 7646
rect 43710 7698 43762 7710
rect 43710 7634 43762 7646
rect 46734 7698 46786 7710
rect 46734 7634 46786 7646
rect 47070 7698 47122 7710
rect 47070 7634 47122 7646
rect 53342 7698 53394 7710
rect 53342 7634 53394 7646
rect 18510 7586 18562 7598
rect 23550 7586 23602 7598
rect 36094 7586 36146 7598
rect 6066 7534 6078 7586
rect 6130 7534 6142 7586
rect 10994 7534 11006 7586
rect 11058 7534 11070 7586
rect 20402 7534 20414 7586
rect 20466 7534 20478 7586
rect 28690 7534 28702 7586
rect 28754 7534 28766 7586
rect 18510 7522 18562 7534
rect 23550 7522 23602 7534
rect 36094 7522 36146 7534
rect 36318 7586 36370 7598
rect 36318 7522 36370 7534
rect 37886 7586 37938 7598
rect 37886 7522 37938 7534
rect 38222 7586 38274 7598
rect 38222 7522 38274 7534
rect 38334 7586 38386 7598
rect 38334 7522 38386 7534
rect 38670 7586 38722 7598
rect 39554 7534 39566 7586
rect 39618 7534 39630 7586
rect 42466 7534 42478 7586
rect 42530 7534 42542 7586
rect 52322 7534 52334 7586
rect 52386 7534 52398 7586
rect 38670 7522 38722 7534
rect 18734 7474 18786 7486
rect 22990 7474 23042 7486
rect 5394 7422 5406 7474
rect 5458 7422 5470 7474
rect 10210 7422 10222 7474
rect 10274 7422 10286 7474
rect 19618 7422 19630 7474
rect 19682 7422 19694 7474
rect 18734 7410 18786 7422
rect 22990 7410 23042 7422
rect 23214 7474 23266 7486
rect 23214 7410 23266 7422
rect 26238 7474 26290 7486
rect 36654 7474 36706 7486
rect 29474 7422 29486 7474
rect 29538 7422 29550 7474
rect 26238 7410 26290 7422
rect 36654 7410 36706 7422
rect 36990 7474 37042 7486
rect 36990 7410 37042 7422
rect 37998 7474 38050 7486
rect 37998 7410 38050 7422
rect 38894 7474 38946 7486
rect 38894 7410 38946 7422
rect 39342 7474 39394 7486
rect 41246 7474 41298 7486
rect 39778 7422 39790 7474
rect 39842 7422 39854 7474
rect 39342 7410 39394 7422
rect 41246 7410 41298 7422
rect 41694 7474 41746 7486
rect 41694 7410 41746 7422
rect 46846 7474 46898 7486
rect 46846 7410 46898 7422
rect 47742 7474 47794 7486
rect 47742 7410 47794 7422
rect 47966 7474 48018 7486
rect 52670 7474 52722 7486
rect 50082 7422 50094 7474
rect 50146 7422 50158 7474
rect 47966 7410 48018 7422
rect 52670 7410 52722 7422
rect 3502 7362 3554 7374
rect 8542 7362 8594 7374
rect 13582 7362 13634 7374
rect 8194 7310 8206 7362
rect 8258 7310 8270 7362
rect 13122 7310 13134 7362
rect 13186 7310 13198 7362
rect 3502 7298 3554 7310
rect 8542 7298 8594 7310
rect 13582 7298 13634 7310
rect 16606 7362 16658 7374
rect 16606 7298 16658 7310
rect 19294 7362 19346 7374
rect 25454 7362 25506 7374
rect 31054 7362 31106 7374
rect 22530 7310 22542 7362
rect 22594 7310 22606 7362
rect 26562 7310 26574 7362
rect 26626 7310 26638 7362
rect 19294 7298 19346 7310
rect 25454 7298 25506 7310
rect 31054 7298 31106 7310
rect 36766 7362 36818 7374
rect 36766 7298 36818 7310
rect 43038 7362 43090 7374
rect 43038 7298 43090 7310
rect 49422 7362 49474 7374
rect 50194 7310 50206 7362
rect 50258 7310 50270 7362
rect 49422 7298 49474 7310
rect 3614 7250 3666 7262
rect 3614 7186 3666 7198
rect 8654 7250 8706 7262
rect 18398 7250 18450 7262
rect 8866 7198 8878 7250
rect 8930 7247 8942 7250
rect 9090 7247 9102 7250
rect 8930 7201 9102 7247
rect 8930 7198 8942 7201
rect 9090 7198 9102 7201
rect 9154 7198 9166 7250
rect 8654 7186 8706 7198
rect 18398 7186 18450 7198
rect 30942 7250 30994 7262
rect 30942 7186 30994 7198
rect 41022 7250 41074 7262
rect 41022 7186 41074 7198
rect 41806 7250 41858 7262
rect 41806 7186 41858 7198
rect 46734 7250 46786 7262
rect 46734 7186 46786 7198
rect 47518 7250 47570 7262
rect 47518 7186 47570 7198
rect 1344 7082 53648 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 53648 7082
rect 1344 6996 53648 7030
rect 32846 6914 32898 6926
rect 32846 6850 32898 6862
rect 39230 6914 39282 6926
rect 39230 6850 39282 6862
rect 43822 6914 43874 6926
rect 43822 6850 43874 6862
rect 49982 6914 50034 6926
rect 49982 6850 50034 6862
rect 48526 6802 48578 6814
rect 16370 6750 16382 6802
rect 16434 6750 16446 6802
rect 19842 6750 19854 6802
rect 19906 6750 19918 6802
rect 45378 6750 45390 6802
rect 45442 6750 45454 6802
rect 48526 6738 48578 6750
rect 8430 6690 8482 6702
rect 8430 6626 8482 6638
rect 8878 6690 8930 6702
rect 9662 6690 9714 6702
rect 27022 6690 27074 6702
rect 9426 6638 9438 6690
rect 9490 6638 9502 6690
rect 13458 6638 13470 6690
rect 13522 6638 13534 6690
rect 14242 6638 14254 6690
rect 14306 6638 14318 6690
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 17714 6638 17726 6690
rect 17778 6638 17790 6690
rect 8878 6626 8930 6638
rect 9662 6626 9714 6638
rect 27022 6626 27074 6638
rect 30718 6690 30770 6702
rect 39118 6690 39170 6702
rect 33506 6638 33518 6690
rect 33570 6638 33582 6690
rect 30718 6626 30770 6638
rect 39118 6626 39170 6638
rect 40798 6690 40850 6702
rect 44046 6690 44098 6702
rect 43362 6638 43374 6690
rect 43426 6638 43438 6690
rect 43586 6638 43598 6690
rect 43650 6638 43662 6690
rect 40798 6626 40850 6638
rect 44046 6626 44098 6638
rect 44830 6690 44882 6702
rect 47630 6690 47682 6702
rect 45714 6638 45726 6690
rect 45778 6638 45790 6690
rect 46498 6638 46510 6690
rect 46562 6638 46574 6690
rect 47394 6638 47406 6690
rect 47458 6638 47470 6690
rect 44830 6626 44882 6638
rect 47630 6626 47682 6638
rect 47854 6690 47906 6702
rect 47854 6626 47906 6638
rect 48078 6690 48130 6702
rect 48078 6626 48130 6638
rect 48414 6690 48466 6702
rect 50206 6690 50258 6702
rect 49746 6638 49758 6690
rect 49810 6638 49822 6690
rect 48414 6626 48466 6638
rect 50206 6626 50258 6638
rect 50430 6690 50482 6702
rect 50430 6626 50482 6638
rect 52670 6690 52722 6702
rect 52670 6626 52722 6638
rect 9998 6578 10050 6590
rect 40910 6578 40962 6590
rect 23874 6526 23886 6578
rect 23938 6526 23950 6578
rect 31378 6526 31390 6578
rect 31442 6526 31454 6578
rect 33394 6526 33406 6578
rect 33458 6526 33470 6578
rect 9998 6514 10050 6526
rect 40910 6514 40962 6526
rect 44270 6578 44322 6590
rect 47182 6578 47234 6590
rect 46274 6526 46286 6578
rect 46338 6526 46350 6578
rect 44270 6514 44322 6526
rect 47182 6514 47234 6526
rect 48862 6578 48914 6590
rect 48862 6514 48914 6526
rect 49534 6578 49586 6590
rect 49534 6514 49586 6526
rect 50766 6578 50818 6590
rect 50766 6514 50818 6526
rect 8990 6466 9042 6478
rect 8990 6402 9042 6414
rect 9102 6466 9154 6478
rect 9102 6402 9154 6414
rect 9886 6466 9938 6478
rect 9886 6402 9938 6414
rect 10558 6466 10610 6478
rect 10558 6402 10610 6414
rect 24222 6466 24274 6478
rect 30382 6466 30434 6478
rect 26674 6414 26686 6466
rect 26738 6414 26750 6466
rect 24222 6402 24274 6414
rect 30382 6402 30434 6414
rect 31054 6466 31106 6478
rect 31054 6402 31106 6414
rect 32510 6466 32562 6478
rect 32510 6402 32562 6414
rect 34190 6466 34242 6478
rect 34190 6402 34242 6414
rect 39230 6466 39282 6478
rect 39230 6402 39282 6414
rect 41134 6466 41186 6478
rect 41134 6402 41186 6414
rect 44382 6466 44434 6478
rect 44382 6402 44434 6414
rect 47630 6466 47682 6478
rect 47630 6402 47682 6414
rect 48638 6466 48690 6478
rect 48638 6402 48690 6414
rect 50542 6466 50594 6478
rect 50542 6402 50594 6414
rect 50878 6466 50930 6478
rect 50878 6402 50930 6414
rect 52222 6466 52274 6478
rect 52222 6402 52274 6414
rect 53230 6466 53282 6478
rect 53230 6402 53282 6414
rect 1344 6298 53648 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 53648 6298
rect 1344 6212 53648 6246
rect 9662 6130 9714 6142
rect 9662 6066 9714 6078
rect 10334 6130 10386 6142
rect 10334 6066 10386 6078
rect 14702 6130 14754 6142
rect 14702 6066 14754 6078
rect 16606 6130 16658 6142
rect 16606 6066 16658 6078
rect 22318 6130 22370 6142
rect 22318 6066 22370 6078
rect 24110 6130 24162 6142
rect 24110 6066 24162 6078
rect 24222 6130 24274 6142
rect 24222 6066 24274 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 27470 6130 27522 6142
rect 27470 6066 27522 6078
rect 27806 6130 27858 6142
rect 27806 6066 27858 6078
rect 9550 6018 9602 6030
rect 9550 5954 9602 5966
rect 14814 6018 14866 6030
rect 14814 5954 14866 5966
rect 22542 6018 22594 6030
rect 22542 5954 22594 5966
rect 22766 6018 22818 6030
rect 34738 5966 34750 6018
rect 34802 5966 34814 6018
rect 51090 5966 51102 6018
rect 51154 5966 51166 6018
rect 22766 5954 22818 5966
rect 22206 5906 22258 5918
rect 22206 5842 22258 5854
rect 24558 5906 24610 5918
rect 24558 5842 24610 5854
rect 27358 5906 27410 5918
rect 27358 5842 27410 5854
rect 27694 5906 27746 5918
rect 48750 5906 48802 5918
rect 33954 5854 33966 5906
rect 34018 5854 34030 5906
rect 49186 5854 49198 5906
rect 49250 5854 49262 5906
rect 50306 5854 50318 5906
rect 50370 5854 50382 5906
rect 27694 5842 27746 5854
rect 48750 5842 48802 5854
rect 22430 5794 22482 5806
rect 22430 5730 22482 5742
rect 24334 5794 24386 5806
rect 24334 5730 24386 5742
rect 27582 5794 27634 5806
rect 37326 5794 37378 5806
rect 36866 5742 36878 5794
rect 36930 5742 36942 5794
rect 27582 5730 27634 5742
rect 37326 5730 37378 5742
rect 49982 5794 50034 5806
rect 53218 5742 53230 5794
rect 53282 5742 53294 5794
rect 49982 5730 50034 5742
rect 9662 5682 9714 5694
rect 9662 5618 9714 5630
rect 1344 5514 53648 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 53648 5514
rect 1344 5428 53648 5462
rect 19518 5346 19570 5358
rect 19518 5282 19570 5294
rect 25006 5346 25058 5358
rect 25006 5282 25058 5294
rect 25342 5346 25394 5358
rect 25342 5282 25394 5294
rect 28142 5346 28194 5358
rect 28142 5282 28194 5294
rect 12350 5234 12402 5246
rect 9762 5182 9774 5234
rect 9826 5182 9838 5234
rect 11890 5182 11902 5234
rect 11954 5182 11966 5234
rect 12350 5170 12402 5182
rect 15598 5234 15650 5246
rect 44942 5234 44994 5246
rect 18834 5182 18846 5234
rect 18898 5182 18910 5234
rect 19170 5182 19182 5234
rect 19234 5182 19246 5234
rect 21298 5182 21310 5234
rect 21362 5182 21374 5234
rect 22418 5182 22430 5234
rect 22482 5182 22494 5234
rect 34066 5182 34078 5234
rect 34130 5182 34142 5234
rect 38770 5182 38782 5234
rect 38834 5182 38846 5234
rect 40898 5182 40910 5234
rect 40962 5182 40974 5234
rect 49522 5182 49534 5234
rect 49586 5182 49598 5234
rect 15598 5170 15650 5182
rect 44942 5170 44994 5182
rect 21646 5122 21698 5134
rect 22542 5122 22594 5134
rect 8978 5070 8990 5122
rect 9042 5070 9054 5122
rect 16034 5070 16046 5122
rect 16098 5070 16110 5122
rect 16706 5070 16718 5122
rect 16770 5070 16782 5122
rect 22306 5070 22318 5122
rect 22370 5070 22382 5122
rect 21646 5058 21698 5070
rect 22542 5058 22594 5070
rect 22766 5122 22818 5134
rect 25790 5122 25842 5134
rect 22978 5070 22990 5122
rect 23042 5070 23054 5122
rect 25330 5070 25342 5122
rect 25394 5070 25406 5122
rect 22766 5058 22818 5070
rect 25790 5058 25842 5070
rect 27806 5122 27858 5134
rect 49982 5122 50034 5134
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 31154 5070 31166 5122
rect 31218 5070 31230 5122
rect 37986 5070 37998 5122
rect 38050 5070 38062 5122
rect 46722 5070 46734 5122
rect 46786 5070 46798 5122
rect 27806 5058 27858 5070
rect 49982 5058 50034 5070
rect 31938 4958 31950 5010
rect 32002 4958 32014 5010
rect 47394 4958 47406 5010
rect 47458 4958 47470 5010
rect 19294 4898 19346 4910
rect 19294 4834 19346 4846
rect 21422 4898 21474 4910
rect 21422 4834 21474 4846
rect 28254 4898 28306 4910
rect 28254 4834 28306 4846
rect 41358 4898 41410 4910
rect 41358 4834 41410 4846
rect 44830 4898 44882 4910
rect 44830 4834 44882 4846
rect 1344 4730 53648 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 53648 4730
rect 1344 4644 53648 4678
rect 14926 4562 14978 4574
rect 14926 4498 14978 4510
rect 31950 4562 32002 4574
rect 31950 4498 32002 4510
rect 44494 4562 44546 4574
rect 44494 4498 44546 4510
rect 47518 4562 47570 4574
rect 47518 4498 47570 4510
rect 48862 4562 48914 4574
rect 48862 4498 48914 4510
rect 49422 4562 49474 4574
rect 49422 4498 49474 4510
rect 25342 4450 25394 4462
rect 32286 4450 32338 4462
rect 47630 4450 47682 4462
rect 20738 4398 20750 4450
rect 20802 4398 20814 4450
rect 29922 4398 29934 4450
rect 29986 4398 29998 4450
rect 36194 4398 36206 4450
rect 36258 4398 36270 4450
rect 41906 4398 41918 4450
rect 41970 4398 41982 4450
rect 25342 4386 25394 4398
rect 32286 4386 32338 4398
rect 47630 4386 47682 4398
rect 49646 4450 49698 4462
rect 49646 4386 49698 4398
rect 49982 4450 50034 4462
rect 51090 4398 51102 4450
rect 51154 4398 51166 4450
rect 49982 4386 50034 4398
rect 19630 4338 19682 4350
rect 38782 4338 38834 4350
rect 14354 4286 14366 4338
rect 14418 4286 14430 4338
rect 19954 4286 19966 4338
rect 20018 4286 20030 4338
rect 30594 4286 30606 4338
rect 30658 4286 30670 4338
rect 35410 4286 35422 4338
rect 35474 4286 35486 4338
rect 41234 4286 41246 4338
rect 41298 4286 41310 4338
rect 50306 4286 50318 4338
rect 50370 4286 50382 4338
rect 19630 4274 19682 4286
rect 38782 4274 38834 4286
rect 48078 4226 48130 4238
rect 22866 4174 22878 4226
rect 22930 4174 22942 4226
rect 27794 4174 27806 4226
rect 27858 4174 27870 4226
rect 38322 4174 38334 4226
rect 38386 4174 38398 4226
rect 44034 4174 44046 4226
rect 44098 4174 44110 4226
rect 53218 4174 53230 4226
rect 53282 4174 53294 4226
rect 48078 4162 48130 4174
rect 12126 4114 12178 4126
rect 12126 4050 12178 4062
rect 1344 3946 53648 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 53648 3946
rect 1344 3860 53648 3894
rect 29822 3666 29874 3678
rect 25330 3614 25342 3666
rect 25394 3614 25406 3666
rect 27458 3614 27470 3666
rect 27522 3614 27534 3666
rect 29822 3602 29874 3614
rect 36990 3666 37042 3678
rect 42030 3666 42082 3678
rect 49646 3666 49698 3678
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 44370 3614 44382 3666
rect 44434 3614 44446 3666
rect 46498 3614 46510 3666
rect 46562 3614 46574 3666
rect 36990 3602 37042 3614
rect 42030 3602 42082 3614
rect 49646 3602 49698 3614
rect 52670 3666 52722 3678
rect 52670 3602 52722 3614
rect 35534 3554 35586 3566
rect 47742 3554 47794 3566
rect 11890 3502 11902 3554
rect 11954 3502 11966 3554
rect 24658 3502 24670 3554
rect 24722 3502 24734 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 50642 3502 50654 3554
rect 50706 3502 50718 3554
rect 35534 3490 35586 3502
rect 47742 3490 47794 3502
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 2942 3442 2994 3454
rect 2942 3378 2994 3390
rect 3278 3442 3330 3454
rect 12462 3442 12514 3454
rect 10098 3390 10110 3442
rect 10162 3390 10174 3442
rect 3278 3378 3330 3390
rect 12462 3378 12514 3390
rect 39342 3442 39394 3454
rect 39342 3378 39394 3390
rect 39790 3442 39842 3454
rect 39790 3378 39842 3390
rect 42478 3442 42530 3454
rect 42478 3378 42530 3390
rect 42702 3442 42754 3454
rect 52446 3442 52498 3454
rect 43026 3390 43038 3442
rect 43090 3390 43102 3442
rect 47394 3390 47406 3442
rect 47458 3390 47470 3442
rect 42702 3378 42754 3390
rect 52446 3378 52498 3390
rect 53230 3442 53282 3454
rect 53230 3378 53282 3390
rect 16942 3330 16994 3342
rect 16942 3266 16994 3278
rect 20862 3330 20914 3342
rect 20862 3266 20914 3278
rect 1344 3162 53648 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 53648 3162
rect 1344 3076 53648 3110
<< via1 >>
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 41246 51550 41298 51602
rect 41470 51550 41522 51602
rect 51214 51326 51266 51378
rect 51438 51326 51490 51378
rect 51662 51326 51714 51378
rect 32398 51214 32450 51266
rect 41918 51214 41970 51266
rect 51326 51214 51378 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 51102 50766 51154 50818
rect 19742 50654 19794 50706
rect 23102 50654 23154 50706
rect 26350 50654 26402 50706
rect 29150 50654 29202 50706
rect 31278 50654 31330 50706
rect 35310 50654 35362 50706
rect 36990 50654 37042 50706
rect 40238 50654 40290 50706
rect 48638 50654 48690 50706
rect 16942 50542 16994 50594
rect 20190 50542 20242 50594
rect 21198 50542 21250 50594
rect 21534 50542 21586 50594
rect 24334 50542 24386 50594
rect 26126 50542 26178 50594
rect 26462 50542 26514 50594
rect 32062 50542 32114 50594
rect 32398 50542 32450 50594
rect 35758 50542 35810 50594
rect 39902 50542 39954 50594
rect 43038 50542 43090 50594
rect 45726 50542 45778 50594
rect 51998 50542 52050 50594
rect 17614 50430 17666 50482
rect 21422 50430 21474 50482
rect 21870 50430 21922 50482
rect 22990 50430 23042 50482
rect 23214 50430 23266 50482
rect 23998 50430 24050 50482
rect 24110 50430 24162 50482
rect 26798 50430 26850 50482
rect 33182 50430 33234 50482
rect 39118 50430 39170 50482
rect 42366 50430 42418 50482
rect 46510 50430 46562 50482
rect 22766 50318 22818 50370
rect 23550 50318 23602 50370
rect 49198 50318 49250 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 20526 49982 20578 50034
rect 21198 49982 21250 50034
rect 21870 49982 21922 50034
rect 26238 49982 26290 50034
rect 33966 49982 34018 50034
rect 36766 49982 36818 50034
rect 37662 49982 37714 50034
rect 41022 49982 41074 50034
rect 49758 49982 49810 50034
rect 49870 49982 49922 50034
rect 49982 49982 50034 50034
rect 21982 49870 22034 49922
rect 23326 49870 23378 49922
rect 23550 49870 23602 49922
rect 25902 49870 25954 49922
rect 26014 49870 26066 49922
rect 27358 49870 27410 49922
rect 27470 49870 27522 49922
rect 33854 49870 33906 49922
rect 37214 49870 37266 49922
rect 37774 49870 37826 49922
rect 41134 49870 41186 49922
rect 43486 49870 43538 49922
rect 48974 49870 49026 49922
rect 51102 49870 51154 49922
rect 19630 49758 19682 49810
rect 19854 49758 19906 49810
rect 21310 49758 21362 49810
rect 26462 49758 26514 49810
rect 26798 49758 26850 49810
rect 26910 49758 26962 49810
rect 27694 49758 27746 49810
rect 32062 49758 32114 49810
rect 33182 49758 33234 49810
rect 34414 49758 34466 49810
rect 34638 49758 34690 49810
rect 34862 49758 34914 49810
rect 35086 49758 35138 49810
rect 36654 49758 36706 49810
rect 36990 49758 37042 49810
rect 39566 49758 39618 49810
rect 39790 49758 39842 49810
rect 40014 49758 40066 49810
rect 40238 49758 40290 49810
rect 42030 49758 42082 49810
rect 42254 49758 42306 49810
rect 42702 49758 42754 49810
rect 48862 49758 48914 49810
rect 49422 49758 49474 49810
rect 50430 49758 50482 49810
rect 23214 49646 23266 49698
rect 26574 49646 26626 49698
rect 28030 49646 28082 49698
rect 29262 49646 29314 49698
rect 31390 49646 31442 49698
rect 34526 49646 34578 49698
rect 36878 49646 36930 49698
rect 37550 49646 37602 49698
rect 39902 49646 39954 49698
rect 40910 49646 40962 49698
rect 45614 49646 45666 49698
rect 53230 49646 53282 49698
rect 20078 49534 20130 49586
rect 21198 49534 21250 49586
rect 21758 49534 21810 49586
rect 34078 49534 34130 49586
rect 42366 49534 42418 49586
rect 48974 49534 49026 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 48750 49198 48802 49250
rect 22094 49086 22146 49138
rect 25678 49086 25730 49138
rect 26462 49086 26514 49138
rect 51886 49086 51938 49138
rect 20750 48974 20802 49026
rect 21646 48974 21698 49026
rect 21758 48974 21810 49026
rect 21982 48974 22034 49026
rect 22654 48974 22706 49026
rect 22990 48974 23042 49026
rect 23438 48974 23490 49026
rect 23662 48974 23714 49026
rect 23998 48974 24050 49026
rect 25566 48974 25618 49026
rect 25790 48974 25842 49026
rect 26014 48974 26066 49026
rect 26350 48974 26402 49026
rect 42702 48974 42754 49026
rect 46062 48974 46114 49026
rect 48974 48974 49026 49026
rect 49198 48974 49250 49026
rect 49646 48974 49698 49026
rect 20414 48862 20466 48914
rect 22430 48862 22482 48914
rect 24558 48862 24610 48914
rect 25342 48862 25394 48914
rect 27134 48862 27186 48914
rect 42254 48862 42306 48914
rect 22766 48750 22818 48802
rect 22878 48750 22930 48802
rect 23550 48750 23602 48802
rect 26574 48750 26626 48802
rect 42478 48750 42530 48802
rect 45950 48750 46002 48802
rect 46398 48750 46450 48802
rect 46622 48750 46674 48802
rect 46734 48750 46786 48802
rect 48302 48750 48354 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 25902 48414 25954 48466
rect 34526 48414 34578 48466
rect 34862 48414 34914 48466
rect 39006 48414 39058 48466
rect 46622 48414 46674 48466
rect 49646 48414 49698 48466
rect 46846 48302 46898 48354
rect 47182 48302 47234 48354
rect 34638 48190 34690 48242
rect 34974 48190 35026 48242
rect 39230 48190 39282 48242
rect 46286 48190 46338 48242
rect 46622 48190 46674 48242
rect 48974 48190 49026 48242
rect 50878 48190 50930 48242
rect 25790 48078 25842 48130
rect 26350 48078 26402 48130
rect 34526 48078 34578 48130
rect 45950 48078 46002 48130
rect 48190 48078 48242 48130
rect 48750 48078 48802 48130
rect 49198 48078 49250 48130
rect 47406 47966 47458 48018
rect 47742 47966 47794 48018
rect 53006 47966 53058 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 27918 47630 27970 47682
rect 37774 47630 37826 47682
rect 12574 47518 12626 47570
rect 19070 47518 19122 47570
rect 34750 47518 34802 47570
rect 42478 47518 42530 47570
rect 49646 47518 49698 47570
rect 51102 47518 51154 47570
rect 9774 47406 9826 47458
rect 16270 47406 16322 47458
rect 20526 47406 20578 47458
rect 20862 47406 20914 47458
rect 21198 47406 21250 47458
rect 21534 47406 21586 47458
rect 28254 47406 28306 47458
rect 31950 47406 32002 47458
rect 39230 47406 39282 47458
rect 42366 47406 42418 47458
rect 42590 47406 42642 47458
rect 42926 47406 42978 47458
rect 49086 47406 49138 47458
rect 49534 47406 49586 47458
rect 10446 47294 10498 47346
rect 16942 47294 16994 47346
rect 20302 47294 20354 47346
rect 21422 47294 21474 47346
rect 21870 47294 21922 47346
rect 24446 47294 24498 47346
rect 24782 47294 24834 47346
rect 25902 47294 25954 47346
rect 32622 47294 32674 47346
rect 35198 47294 35250 47346
rect 36990 47294 37042 47346
rect 37662 47294 37714 47346
rect 37774 47294 37826 47346
rect 38334 47294 38386 47346
rect 39454 47294 39506 47346
rect 48750 47294 48802 47346
rect 50430 47294 50482 47346
rect 50766 47294 50818 47346
rect 9326 47182 9378 47234
rect 19406 47182 19458 47234
rect 19742 47182 19794 47234
rect 20750 47182 20802 47234
rect 26238 47182 26290 47234
rect 28030 47182 28082 47234
rect 31166 47182 31218 47234
rect 31502 47182 31554 47234
rect 37326 47182 37378 47234
rect 42814 47182 42866 47234
rect 46846 47182 46898 47234
rect 48862 47182 48914 47234
rect 50990 47182 51042 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 17950 46846 18002 46898
rect 19294 46846 19346 46898
rect 20974 46846 21026 46898
rect 24110 46846 24162 46898
rect 33182 46846 33234 46898
rect 37102 46846 37154 46898
rect 41806 46846 41858 46898
rect 42142 46846 42194 46898
rect 20526 46734 20578 46786
rect 21086 46734 21138 46786
rect 30046 46734 30098 46786
rect 33406 46734 33458 46786
rect 41582 46734 41634 46786
rect 42926 46734 42978 46786
rect 47854 46734 47906 46786
rect 51102 46734 51154 46786
rect 13022 46622 13074 46674
rect 16158 46622 16210 46674
rect 16382 46622 16434 46674
rect 16606 46622 16658 46674
rect 17502 46622 17554 46674
rect 20638 46622 20690 46674
rect 23102 46622 23154 46674
rect 23214 46622 23266 46674
rect 23326 46622 23378 46674
rect 23774 46622 23826 46674
rect 26238 46622 26290 46674
rect 30718 46622 30770 46674
rect 36430 46622 36482 46674
rect 36878 46622 36930 46674
rect 37438 46622 37490 46674
rect 41246 46622 41298 46674
rect 42030 46622 42082 46674
rect 43374 46622 43426 46674
rect 47742 46622 47794 46674
rect 48078 46622 48130 46674
rect 50430 46622 50482 46674
rect 13694 46510 13746 46562
rect 15822 46510 15874 46562
rect 16270 46510 16322 46562
rect 26798 46510 26850 46562
rect 27918 46510 27970 46562
rect 31166 46510 31218 46562
rect 31278 46510 31330 46562
rect 17390 46398 17442 46450
rect 20526 46398 20578 46450
rect 31726 46510 31778 46562
rect 33070 46510 33122 46562
rect 36206 46510 36258 46562
rect 36990 46510 37042 46562
rect 38222 46510 38274 46562
rect 40350 46510 40402 46562
rect 41918 46510 41970 46562
rect 43038 46510 43090 46562
rect 44158 46510 44210 46562
rect 46286 46510 46338 46562
rect 53230 46510 53282 46562
rect 31838 46398 31890 46450
rect 42702 46398 42754 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 16270 46062 16322 46114
rect 21646 46062 21698 46114
rect 10894 45950 10946 46002
rect 34750 45950 34802 46002
rect 37998 45950 38050 46002
rect 42702 45950 42754 46002
rect 45390 45950 45442 46002
rect 48078 45950 48130 46002
rect 10782 45838 10834 45890
rect 11118 45838 11170 45890
rect 16382 45838 16434 45890
rect 16830 45838 16882 45890
rect 16942 45838 16994 45890
rect 17390 45838 17442 45890
rect 21982 45838 22034 45890
rect 22206 45838 22258 45890
rect 22654 45838 22706 45890
rect 22766 45838 22818 45890
rect 25902 45838 25954 45890
rect 36990 45838 37042 45890
rect 37550 45838 37602 45890
rect 42590 45838 42642 45890
rect 42814 45838 42866 45890
rect 43038 45838 43090 45890
rect 47070 45838 47122 45890
rect 48190 45838 48242 45890
rect 49198 45838 49250 45890
rect 49422 45838 49474 45890
rect 10446 45726 10498 45778
rect 11454 45726 11506 45778
rect 17614 45726 17666 45778
rect 17950 45726 18002 45778
rect 18510 45726 18562 45778
rect 24110 45726 24162 45778
rect 25342 45726 25394 45778
rect 25790 45726 25842 45778
rect 26014 45726 26066 45778
rect 26238 45726 26290 45778
rect 35086 45726 35138 45778
rect 37214 45726 37266 45778
rect 42366 45726 42418 45778
rect 47742 45726 47794 45778
rect 49086 45726 49138 45778
rect 15934 45614 15986 45666
rect 16270 45614 16322 45666
rect 16718 45614 16770 45666
rect 22878 45614 22930 45666
rect 22990 45614 23042 45666
rect 23102 45614 23154 45666
rect 24446 45614 24498 45666
rect 25118 45614 25170 45666
rect 26350 45614 26402 45666
rect 34862 45614 34914 45666
rect 37438 45614 37490 45666
rect 44270 45614 44322 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 11006 45278 11058 45330
rect 14814 45278 14866 45330
rect 17502 45278 17554 45330
rect 23102 45278 23154 45330
rect 23214 45278 23266 45330
rect 24670 45278 24722 45330
rect 41246 45278 41298 45330
rect 41918 45278 41970 45330
rect 48078 45278 48130 45330
rect 48750 45278 48802 45330
rect 12238 45166 12290 45218
rect 12910 45166 12962 45218
rect 19966 45166 20018 45218
rect 28814 45166 28866 45218
rect 33070 45166 33122 45218
rect 38334 45166 38386 45218
rect 38894 45166 38946 45218
rect 42254 45166 42306 45218
rect 42478 45166 42530 45218
rect 43710 45166 43762 45218
rect 48190 45166 48242 45218
rect 48862 45166 48914 45218
rect 10894 45054 10946 45106
rect 11118 45054 11170 45106
rect 11566 45054 11618 45106
rect 11790 45054 11842 45106
rect 12014 45054 12066 45106
rect 12462 45054 12514 45106
rect 13358 45054 13410 45106
rect 13918 45054 13970 45106
rect 14254 45054 14306 45106
rect 17278 45054 17330 45106
rect 17614 45054 17666 45106
rect 18734 45054 18786 45106
rect 19518 45054 19570 45106
rect 20078 45054 20130 45106
rect 21870 45054 21922 45106
rect 22094 45054 22146 45106
rect 25678 45054 25730 45106
rect 29038 45054 29090 45106
rect 29598 45054 29650 45106
rect 31950 45054 32002 45106
rect 32398 45054 32450 45106
rect 33630 45054 33682 45106
rect 34190 45054 34242 45106
rect 37214 45054 37266 45106
rect 38222 45054 38274 45106
rect 41134 45054 41186 45106
rect 46622 45054 46674 45106
rect 47854 45054 47906 45106
rect 50318 45054 50370 45106
rect 12910 44942 12962 44994
rect 14366 44942 14418 44994
rect 22430 44942 22482 44994
rect 22990 44942 23042 44994
rect 26350 44942 26402 44994
rect 28478 44942 28530 44994
rect 31614 44942 31666 44994
rect 33854 44942 33906 44994
rect 34862 44942 34914 44994
rect 35646 44942 35698 44994
rect 39454 44942 39506 44994
rect 42366 44942 42418 44994
rect 45278 44942 45330 44994
rect 47518 44942 47570 44994
rect 49982 44942 50034 44994
rect 51102 44942 51154 44994
rect 53230 44942 53282 44994
rect 12350 44830 12402 44882
rect 19854 44830 19906 44882
rect 22318 44830 22370 44882
rect 41246 44830 41298 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 25902 44494 25954 44546
rect 26238 44494 26290 44546
rect 33294 44494 33346 44546
rect 35534 44494 35586 44546
rect 38446 44494 38498 44546
rect 38894 44494 38946 44546
rect 9662 44382 9714 44434
rect 10110 44382 10162 44434
rect 22094 44382 22146 44434
rect 32062 44382 32114 44434
rect 35086 44382 35138 44434
rect 39454 44382 39506 44434
rect 42142 44382 42194 44434
rect 44270 44382 44322 44434
rect 51774 44382 51826 44434
rect 6862 44270 6914 44322
rect 10670 44270 10722 44322
rect 11342 44270 11394 44322
rect 11790 44270 11842 44322
rect 12574 44270 12626 44322
rect 12686 44270 12738 44322
rect 12798 44270 12850 44322
rect 14478 44270 14530 44322
rect 15934 44270 15986 44322
rect 16494 44270 16546 44322
rect 17278 44270 17330 44322
rect 17502 44270 17554 44322
rect 19294 44270 19346 44322
rect 19742 44270 19794 44322
rect 19966 44270 20018 44322
rect 21310 44270 21362 44322
rect 25118 44270 25170 44322
rect 29262 44270 29314 44322
rect 32398 44270 32450 44322
rect 32622 44270 32674 44322
rect 32846 44270 32898 44322
rect 33630 44270 33682 44322
rect 34078 44270 34130 44322
rect 34750 44270 34802 44322
rect 36094 44270 36146 44322
rect 36318 44270 36370 44322
rect 38558 44270 38610 44322
rect 39006 44270 39058 44322
rect 41358 44270 41410 44322
rect 45054 44270 45106 44322
rect 45614 44270 45666 44322
rect 45950 44270 46002 44322
rect 47518 44270 47570 44322
rect 51102 44270 51154 44322
rect 51214 44270 51266 44322
rect 51662 44270 51714 44322
rect 7534 44158 7586 44210
rect 11678 44158 11730 44210
rect 16046 44158 16098 44210
rect 17838 44158 17890 44210
rect 19854 44158 19906 44210
rect 22542 44158 22594 44210
rect 23998 44158 24050 44210
rect 26126 44158 26178 44210
rect 29934 44158 29986 44210
rect 34414 44158 34466 44210
rect 35758 44158 35810 44210
rect 38222 44158 38274 44210
rect 39790 44158 39842 44210
rect 39902 44158 39954 44210
rect 40686 44158 40738 44210
rect 44942 44158 44994 44210
rect 45502 44158 45554 44210
rect 46062 44158 46114 44210
rect 10782 44046 10834 44098
rect 10894 44046 10946 44098
rect 11454 44046 11506 44098
rect 12126 44046 12178 44098
rect 14702 44046 14754 44098
rect 15150 44046 15202 44098
rect 16158 44046 16210 44098
rect 16830 44046 16882 44098
rect 17390 44046 17442 44098
rect 36430 44046 36482 44098
rect 40126 44046 40178 44098
rect 40350 44046 40402 44098
rect 44718 44046 44770 44098
rect 45278 44046 45330 44098
rect 46286 44046 46338 44098
rect 47742 44046 47794 44098
rect 50878 44046 50930 44098
rect 51326 44046 51378 44098
rect 51886 44046 51938 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 11118 43710 11170 43762
rect 39230 43710 39282 43762
rect 47630 43710 47682 43762
rect 9662 43598 9714 43650
rect 9774 43598 9826 43650
rect 9998 43598 10050 43650
rect 19406 43598 19458 43650
rect 20078 43598 20130 43650
rect 21310 43598 21362 43650
rect 22430 43598 22482 43650
rect 28814 43598 28866 43650
rect 34526 43598 34578 43650
rect 37886 43598 37938 43650
rect 39454 43598 39506 43650
rect 44494 43598 44546 43650
rect 10222 43486 10274 43538
rect 10894 43486 10946 43538
rect 16270 43486 16322 43538
rect 16494 43486 16546 43538
rect 19742 43486 19794 43538
rect 20414 43486 20466 43538
rect 21646 43486 21698 43538
rect 22766 43486 22818 43538
rect 32286 43486 32338 43538
rect 33070 43486 33122 43538
rect 34190 43486 34242 43538
rect 34862 43486 34914 43538
rect 37774 43486 37826 43538
rect 38782 43486 38834 43538
rect 40014 43486 40066 43538
rect 41470 43486 41522 43538
rect 47294 43486 47346 43538
rect 51102 43486 51154 43538
rect 17614 43374 17666 43426
rect 31502 43374 31554 43426
rect 32398 43374 32450 43426
rect 33518 43374 33570 43426
rect 35982 43374 36034 43426
rect 39790 43374 39842 43426
rect 41134 43374 41186 43426
rect 41918 43374 41970 43426
rect 46846 43374 46898 43426
rect 47070 43374 47122 43426
rect 53006 43374 53058 43426
rect 16718 43262 16770 43314
rect 16830 43262 16882 43314
rect 31950 43262 32002 43314
rect 32062 43262 32114 43314
rect 34190 43262 34242 43314
rect 40350 43262 40402 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 23550 42926 23602 42978
rect 33742 42926 33794 42978
rect 34078 42926 34130 42978
rect 34862 42926 34914 42978
rect 15486 42814 15538 42866
rect 17614 42814 17666 42866
rect 18062 42814 18114 42866
rect 25454 42814 25506 42866
rect 26350 42814 26402 42866
rect 26686 42814 26738 42866
rect 32398 42814 32450 42866
rect 32734 42814 32786 42866
rect 33854 42814 33906 42866
rect 46734 42814 46786 42866
rect 47854 42814 47906 42866
rect 49982 42814 50034 42866
rect 50990 42814 51042 42866
rect 12462 42702 12514 42754
rect 14814 42702 14866 42754
rect 19182 42702 19234 42754
rect 23662 42702 23714 42754
rect 23886 42702 23938 42754
rect 24110 42702 24162 42754
rect 25006 42702 25058 42754
rect 27918 42702 27970 42754
rect 28366 42702 28418 42754
rect 29262 42702 29314 42754
rect 29486 42702 29538 42754
rect 29710 42702 29762 42754
rect 38558 42702 38610 42754
rect 40014 42702 40066 42754
rect 47070 42702 47122 42754
rect 19070 42590 19122 42642
rect 24446 42590 24498 42642
rect 25230 42590 25282 42642
rect 25566 42590 25618 42642
rect 26014 42590 26066 42642
rect 26574 42590 26626 42642
rect 35870 42590 35922 42642
rect 35982 42590 36034 42642
rect 39902 42590 39954 42642
rect 50654 42590 50706 42642
rect 50878 42590 50930 42642
rect 10446 42478 10498 42530
rect 10894 42478 10946 42530
rect 12574 42478 12626 42530
rect 12798 42478 12850 42530
rect 18846 42478 18898 42530
rect 24670 42478 24722 42530
rect 24782 42478 24834 42530
rect 27470 42478 27522 42530
rect 28590 42478 28642 42530
rect 29598 42478 29650 42530
rect 34414 42478 34466 42530
rect 34750 42478 34802 42530
rect 36206 42478 36258 42530
rect 38222 42478 38274 42530
rect 39678 42478 39730 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 11678 42142 11730 42194
rect 12686 42142 12738 42194
rect 13246 42142 13298 42194
rect 23886 42142 23938 42194
rect 24670 42142 24722 42194
rect 25566 42142 25618 42194
rect 25790 42142 25842 42194
rect 34414 42142 34466 42194
rect 34974 42142 35026 42194
rect 49758 42142 49810 42194
rect 10894 42030 10946 42082
rect 11118 42030 11170 42082
rect 11230 42030 11282 42082
rect 13022 42030 13074 42082
rect 27022 42030 27074 42082
rect 33406 42030 33458 42082
rect 33518 42030 33570 42082
rect 34526 42030 34578 42082
rect 35086 42030 35138 42082
rect 41246 42030 41298 42082
rect 49982 42030 50034 42082
rect 51102 42030 51154 42082
rect 10222 41918 10274 41970
rect 10446 41918 10498 41970
rect 10782 41918 10834 41970
rect 12350 41918 12402 41970
rect 12910 41918 12962 41970
rect 13470 41918 13522 41970
rect 21982 41918 22034 41970
rect 23102 41918 23154 41970
rect 23214 41918 23266 41970
rect 23662 41918 23714 41970
rect 24222 41918 24274 41970
rect 24558 41918 24610 41970
rect 25118 41918 25170 41970
rect 26350 41918 26402 41970
rect 29822 41918 29874 41970
rect 33742 41918 33794 41970
rect 34190 41918 34242 41970
rect 41022 41918 41074 41970
rect 41694 41918 41746 41970
rect 47406 41918 47458 41970
rect 47966 41918 48018 41970
rect 49086 41918 49138 41970
rect 49310 41918 49362 41970
rect 49870 41918 49922 41970
rect 50318 41918 50370 41970
rect 10558 41806 10610 41858
rect 12126 41806 12178 41858
rect 23438 41806 23490 41858
rect 25678 41806 25730 41858
rect 29150 41806 29202 41858
rect 41470 41806 41522 41858
rect 44606 41806 44658 41858
rect 46734 41806 46786 41858
rect 53230 41806 53282 41858
rect 34974 41694 35026 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14030 41358 14082 41410
rect 22430 41358 22482 41410
rect 8094 41246 8146 41298
rect 10222 41246 10274 41298
rect 14814 41246 14866 41298
rect 20526 41246 20578 41298
rect 26126 41246 26178 41298
rect 33182 41246 33234 41298
rect 38558 41246 38610 41298
rect 40910 41246 40962 41298
rect 43038 41246 43090 41298
rect 43486 41246 43538 41298
rect 48526 41246 48578 41298
rect 51886 41246 51938 41298
rect 7310 41134 7362 41186
rect 10894 41134 10946 41186
rect 12350 41134 12402 41186
rect 12686 41134 12738 41186
rect 13470 41134 13522 41186
rect 13694 41134 13746 41186
rect 14030 41134 14082 41186
rect 17726 41134 17778 41186
rect 18286 41134 18338 41186
rect 18734 41134 18786 41186
rect 18958 41134 19010 41186
rect 19966 41134 20018 41186
rect 20414 41134 20466 41186
rect 20638 41134 20690 41186
rect 21758 41134 21810 41186
rect 22654 41134 22706 41186
rect 22878 41134 22930 41186
rect 30382 41134 30434 41186
rect 33742 41134 33794 41186
rect 34078 41134 34130 41186
rect 37102 41134 37154 41186
rect 37214 41134 37266 41186
rect 38110 41134 38162 41186
rect 39678 41134 39730 41186
rect 40126 41134 40178 41186
rect 44382 41134 44434 41186
rect 44718 41134 44770 41186
rect 45166 41134 45218 41186
rect 48862 41134 48914 41186
rect 49982 41134 50034 41186
rect 11118 41022 11170 41074
rect 12910 41022 12962 41074
rect 18062 41022 18114 41074
rect 18510 41022 18562 41074
rect 19182 41022 19234 41074
rect 20190 41022 20242 41074
rect 21198 41022 21250 41074
rect 21310 41022 21362 41074
rect 31054 41022 31106 41074
rect 33854 41022 33906 41074
rect 34302 41022 34354 41074
rect 37550 41022 37602 41074
rect 37774 41022 37826 41074
rect 44046 41022 44098 41074
rect 45390 41022 45442 41074
rect 49198 41022 49250 41074
rect 11566 40910 11618 40962
rect 13022 40910 13074 40962
rect 13918 40910 13970 40962
rect 17838 40910 17890 40962
rect 18622 40910 18674 40962
rect 19630 40910 19682 40962
rect 21534 40910 21586 40962
rect 22766 40910 22818 40962
rect 37326 40910 37378 40962
rect 37998 40910 38050 40962
rect 39454 40910 39506 40962
rect 44158 40910 44210 40962
rect 45054 40910 45106 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 10782 40574 10834 40626
rect 19182 40574 19234 40626
rect 20526 40574 20578 40626
rect 30046 40574 30098 40626
rect 30382 40574 30434 40626
rect 30718 40574 30770 40626
rect 31390 40574 31442 40626
rect 40910 40574 40962 40626
rect 41694 40574 41746 40626
rect 21758 40462 21810 40514
rect 22430 40462 22482 40514
rect 33966 40462 34018 40514
rect 34190 40462 34242 40514
rect 36654 40462 36706 40514
rect 41246 40462 41298 40514
rect 41918 40462 41970 40514
rect 19070 40350 19122 40402
rect 20302 40350 20354 40402
rect 20862 40350 20914 40402
rect 23998 40350 24050 40402
rect 31054 40350 31106 40402
rect 33854 40350 33906 40402
rect 34302 40350 34354 40402
rect 35870 40350 35922 40402
rect 42030 40350 42082 40402
rect 44942 40350 44994 40402
rect 45278 40350 45330 40402
rect 45502 40350 45554 40402
rect 50654 40350 50706 40402
rect 14590 40238 14642 40290
rect 21870 40238 21922 40290
rect 33406 40238 33458 40290
rect 38782 40238 38834 40290
rect 39230 40238 39282 40290
rect 45166 40238 45218 40290
rect 14254 40126 14306 40178
rect 14590 40126 14642 40178
rect 53006 40126 53058 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 13918 39790 13970 39842
rect 14590 39790 14642 39842
rect 44942 39790 44994 39842
rect 8542 39678 8594 39730
rect 8990 39678 9042 39730
rect 16158 39678 16210 39730
rect 18398 39678 18450 39730
rect 18958 39678 19010 39730
rect 21646 39678 21698 39730
rect 22766 39678 22818 39730
rect 24894 39678 24946 39730
rect 25902 39678 25954 39730
rect 26126 39678 26178 39730
rect 26350 39678 26402 39730
rect 46062 39678 46114 39730
rect 46398 39678 46450 39730
rect 48526 39678 48578 39730
rect 50878 39678 50930 39730
rect 5742 39566 5794 39618
rect 10110 39566 10162 39618
rect 10558 39566 10610 39618
rect 11006 39566 11058 39618
rect 13806 39566 13858 39618
rect 14254 39566 14306 39618
rect 15486 39566 15538 39618
rect 22094 39566 22146 39618
rect 25230 39566 25282 39618
rect 25566 39566 25618 39618
rect 25790 39566 25842 39618
rect 28142 39566 28194 39618
rect 28366 39566 28418 39618
rect 33518 39566 33570 39618
rect 33854 39566 33906 39618
rect 34190 39566 34242 39618
rect 49198 39566 49250 39618
rect 6414 39454 6466 39506
rect 11230 39454 11282 39506
rect 13470 39454 13522 39506
rect 14702 39454 14754 39506
rect 28590 39454 28642 39506
rect 44830 39454 44882 39506
rect 50542 39454 50594 39506
rect 50766 39454 50818 39506
rect 11678 39342 11730 39394
rect 13918 39342 13970 39394
rect 25342 39342 25394 39394
rect 29262 39342 29314 39394
rect 30718 39342 30770 39394
rect 33630 39342 33682 39394
rect 44942 39342 44994 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 6862 39006 6914 39058
rect 10110 39006 10162 39058
rect 10558 39006 10610 39058
rect 15374 39006 15426 39058
rect 17838 39006 17890 39058
rect 24558 39006 24610 39058
rect 29374 39006 29426 39058
rect 33182 39006 33234 39058
rect 41134 39006 41186 39058
rect 44382 39006 44434 39058
rect 49870 39006 49922 39058
rect 49982 39006 50034 39058
rect 9774 38894 9826 38946
rect 12798 38894 12850 38946
rect 18958 38894 19010 38946
rect 29150 38894 29202 38946
rect 30382 38894 30434 38946
rect 40126 38894 40178 38946
rect 40238 38894 40290 38946
rect 41246 38894 41298 38946
rect 44942 38894 44994 38946
rect 45054 38894 45106 38946
rect 51102 38894 51154 38946
rect 6526 38782 6578 38834
rect 6862 38782 6914 38834
rect 7086 38782 7138 38834
rect 12126 38782 12178 38834
rect 18174 38782 18226 38834
rect 23998 38782 24050 38834
rect 27022 38782 27074 38834
rect 27470 38782 27522 38834
rect 29038 38782 29090 38834
rect 29710 38782 29762 38834
rect 35422 38782 35474 38834
rect 40462 38782 40514 38834
rect 40798 38782 40850 38834
rect 41358 38782 41410 38834
rect 44046 38782 44098 38834
rect 44382 38782 44434 38834
rect 44718 38782 44770 38834
rect 49310 38782 49362 38834
rect 49758 38782 49810 38834
rect 50430 38782 50482 38834
rect 14926 38670 14978 38722
rect 21086 38670 21138 38722
rect 27918 38670 27970 38722
rect 28478 38670 28530 38722
rect 32510 38670 32562 38722
rect 36094 38670 36146 38722
rect 38222 38670 38274 38722
rect 38894 38670 38946 38722
rect 53230 38670 53282 38722
rect 45054 38558 45106 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 6862 38222 6914 38274
rect 29150 38222 29202 38274
rect 29710 38222 29762 38274
rect 29822 38222 29874 38274
rect 35982 38110 36034 38162
rect 37102 38110 37154 38162
rect 39230 38110 39282 38162
rect 41358 38110 41410 38162
rect 49982 38110 50034 38162
rect 6974 37998 7026 38050
rect 28142 37998 28194 38050
rect 28366 37998 28418 38050
rect 28590 37998 28642 38050
rect 29262 37998 29314 38050
rect 29486 37998 29538 38050
rect 33070 37998 33122 38050
rect 42142 37998 42194 38050
rect 33742 37886 33794 37938
rect 38110 37886 38162 37938
rect 6862 37774 6914 37826
rect 27246 37774 27298 37826
rect 37774 37774 37826 37826
rect 42590 37774 42642 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 19182 37438 19234 37490
rect 46286 37438 46338 37490
rect 49422 37438 49474 37490
rect 49646 37438 49698 37490
rect 5182 37326 5234 37378
rect 7086 37326 7138 37378
rect 7422 37326 7474 37378
rect 18958 37326 19010 37378
rect 19630 37326 19682 37378
rect 26126 37326 26178 37378
rect 29262 37326 29314 37378
rect 43710 37326 43762 37378
rect 1822 37214 1874 37266
rect 5294 37214 5346 37266
rect 5630 37214 5682 37266
rect 5854 37214 5906 37266
rect 6190 37214 6242 37266
rect 6638 37214 6690 37266
rect 6862 37214 6914 37266
rect 9550 37214 9602 37266
rect 13694 37214 13746 37266
rect 14926 37214 14978 37266
rect 15374 37214 15426 37266
rect 16158 37214 16210 37266
rect 17838 37214 17890 37266
rect 18846 37214 18898 37266
rect 20526 37214 20578 37266
rect 25902 37214 25954 37266
rect 28814 37214 28866 37266
rect 29150 37214 29202 37266
rect 42926 37214 42978 37266
rect 48190 37214 48242 37266
rect 48974 37214 49026 37266
rect 50654 37214 50706 37266
rect 2494 37102 2546 37154
rect 4622 37102 4674 37154
rect 5742 37102 5794 37154
rect 6974 37102 7026 37154
rect 7534 37102 7586 37154
rect 8990 37102 9042 37154
rect 10334 37102 10386 37154
rect 12462 37102 12514 37154
rect 13806 37102 13858 37154
rect 14142 37102 14194 37154
rect 15486 37102 15538 37154
rect 16382 37102 16434 37154
rect 16830 37102 16882 37154
rect 18174 37102 18226 37154
rect 18510 37102 18562 37154
rect 19854 37102 19906 37154
rect 20750 37102 20802 37154
rect 21422 37102 21474 37154
rect 22990 37102 23042 37154
rect 29822 37102 29874 37154
rect 37438 37102 37490 37154
rect 45838 37102 45890 37154
rect 49534 37102 49586 37154
rect 5182 36990 5234 37042
rect 53006 36990 53058 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 5742 36654 5794 36706
rect 9998 36542 10050 36594
rect 17950 36542 18002 36594
rect 23998 36542 24050 36594
rect 25678 36542 25730 36594
rect 45726 36542 45778 36594
rect 47294 36542 47346 36594
rect 49422 36542 49474 36594
rect 5518 36430 5570 36482
rect 15710 36430 15762 36482
rect 17166 36430 17218 36482
rect 18286 36430 18338 36482
rect 22094 36430 22146 36482
rect 22542 36430 22594 36482
rect 23102 36430 23154 36482
rect 23550 36430 23602 36482
rect 24894 36430 24946 36482
rect 25342 36430 25394 36482
rect 39118 36430 39170 36482
rect 39342 36430 39394 36482
rect 40574 36430 40626 36482
rect 43710 36430 43762 36482
rect 44830 36430 44882 36482
rect 45502 36430 45554 36482
rect 46174 36430 46226 36482
rect 46510 36430 46562 36482
rect 50990 36430 51042 36482
rect 51214 36430 51266 36482
rect 9550 36318 9602 36370
rect 10222 36318 10274 36370
rect 16606 36318 16658 36370
rect 18174 36318 18226 36370
rect 22654 36318 22706 36370
rect 24334 36318 24386 36370
rect 26014 36318 26066 36370
rect 40686 36318 40738 36370
rect 42254 36318 42306 36370
rect 42366 36318 42418 36370
rect 43822 36318 43874 36370
rect 44942 36318 44994 36370
rect 45950 36318 46002 36370
rect 4846 36206 4898 36258
rect 5854 36206 5906 36258
rect 6078 36206 6130 36258
rect 9214 36206 9266 36258
rect 9998 36206 10050 36258
rect 10670 36206 10722 36258
rect 38334 36206 38386 36258
rect 38782 36206 38834 36258
rect 38894 36206 38946 36258
rect 39006 36206 39058 36258
rect 40910 36206 40962 36258
rect 42030 36206 42082 36258
rect 42926 36206 42978 36258
rect 44046 36206 44098 36258
rect 45166 36206 45218 36258
rect 50766 36206 50818 36258
rect 51102 36206 51154 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 5294 35870 5346 35922
rect 5742 35870 5794 35922
rect 6862 35870 6914 35922
rect 6974 35870 7026 35922
rect 9998 35870 10050 35922
rect 16606 35870 16658 35922
rect 32622 35870 32674 35922
rect 43038 35870 43090 35922
rect 44158 35870 44210 35922
rect 44382 35870 44434 35922
rect 46174 35870 46226 35922
rect 49982 35870 50034 35922
rect 5182 35758 5234 35810
rect 5406 35758 5458 35810
rect 6302 35758 6354 35810
rect 7310 35758 7362 35810
rect 9550 35758 9602 35810
rect 22878 35758 22930 35810
rect 26238 35758 26290 35810
rect 30606 35758 30658 35810
rect 32398 35758 32450 35810
rect 34078 35758 34130 35810
rect 40910 35758 40962 35810
rect 44830 35758 44882 35810
rect 6190 35646 6242 35698
rect 6526 35646 6578 35698
rect 7086 35646 7138 35698
rect 9774 35646 9826 35698
rect 11790 35646 11842 35698
rect 12126 35646 12178 35698
rect 12910 35646 12962 35698
rect 13358 35646 13410 35698
rect 15598 35646 15650 35698
rect 16046 35646 16098 35698
rect 17838 35646 17890 35698
rect 18286 35646 18338 35698
rect 19294 35646 19346 35698
rect 19742 35646 19794 35698
rect 20414 35646 20466 35698
rect 22206 35646 22258 35698
rect 25790 35646 25842 35698
rect 26798 35646 26850 35698
rect 30158 35646 30210 35698
rect 30942 35646 30994 35698
rect 31614 35646 31666 35698
rect 32174 35646 32226 35698
rect 33182 35646 33234 35698
rect 33966 35646 34018 35698
rect 34302 35646 34354 35698
rect 35422 35646 35474 35698
rect 38894 35646 38946 35698
rect 41134 35646 41186 35698
rect 41694 35646 41746 35698
rect 42142 35646 42194 35698
rect 42702 35646 42754 35698
rect 43710 35646 43762 35698
rect 43934 35646 43986 35698
rect 44382 35646 44434 35698
rect 50318 35646 50370 35698
rect 9998 35534 10050 35586
rect 12238 35534 12290 35586
rect 13582 35534 13634 35586
rect 14030 35534 14082 35586
rect 15150 35534 15202 35586
rect 18510 35534 18562 35586
rect 19854 35534 19906 35586
rect 21982 35534 22034 35586
rect 23438 35534 23490 35586
rect 24222 35534 24274 35586
rect 25342 35534 25394 35586
rect 27134 35534 27186 35586
rect 29038 35534 29090 35586
rect 29486 35534 29538 35586
rect 34638 35534 34690 35586
rect 36094 35534 36146 35586
rect 38222 35534 38274 35586
rect 39790 35534 39842 35586
rect 40350 35534 40402 35586
rect 45278 35534 45330 35586
rect 49198 35534 49250 35586
rect 51102 35534 51154 35586
rect 53230 35534 53282 35586
rect 34414 35422 34466 35474
rect 34862 35422 34914 35474
rect 42478 35422 42530 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 33854 35086 33906 35138
rect 36094 35086 36146 35138
rect 50878 35086 50930 35138
rect 4622 34974 4674 35026
rect 5182 34974 5234 35026
rect 8430 34974 8482 35026
rect 10222 34974 10274 35026
rect 11566 34974 11618 35026
rect 12462 34974 12514 35026
rect 17502 34974 17554 35026
rect 30158 34974 30210 35026
rect 31726 34974 31778 35026
rect 35086 34974 35138 35026
rect 38446 34974 38498 35026
rect 40126 34974 40178 35026
rect 45166 34974 45218 35026
rect 46734 34974 46786 35026
rect 48862 34974 48914 35026
rect 51102 34974 51154 35026
rect 1822 34862 1874 34914
rect 7534 34862 7586 34914
rect 9886 34862 9938 34914
rect 10334 34862 10386 34914
rect 15710 34862 15762 34914
rect 19070 34862 19122 34914
rect 19630 34862 19682 34914
rect 31054 34862 31106 34914
rect 31950 34862 32002 34914
rect 32622 34862 32674 34914
rect 32958 34862 33010 34914
rect 33630 34862 33682 34914
rect 38894 34862 38946 34914
rect 39230 34862 39282 34914
rect 39790 34862 39842 34914
rect 41582 34862 41634 34914
rect 45278 34862 45330 34914
rect 45950 34862 46002 34914
rect 49534 34862 49586 34914
rect 49758 34862 49810 34914
rect 2494 34750 2546 34802
rect 18510 34750 18562 34802
rect 20078 34750 20130 34802
rect 25342 34750 25394 34802
rect 25678 34750 25730 34802
rect 31278 34750 31330 34802
rect 33406 34750 33458 34802
rect 34750 34750 34802 34802
rect 35534 34750 35586 34802
rect 39454 34750 39506 34802
rect 40462 34750 40514 34802
rect 42478 34750 42530 34802
rect 42590 34750 42642 34802
rect 45054 34750 45106 34802
rect 45614 34750 45666 34802
rect 49646 34750 49698 34802
rect 10110 34638 10162 34690
rect 10446 34638 10498 34690
rect 11006 34638 11058 34690
rect 18174 34638 18226 34690
rect 19182 34638 19234 34690
rect 26126 34638 26178 34690
rect 29710 34638 29762 34690
rect 30606 34638 30658 34690
rect 33966 34638 34018 34690
rect 34190 34638 34242 34690
rect 34974 34638 35026 34690
rect 35198 34638 35250 34690
rect 35758 34638 35810 34690
rect 35982 34638 36034 34690
rect 39006 34638 39058 34690
rect 39118 34638 39170 34690
rect 40014 34638 40066 34690
rect 40238 34638 40290 34690
rect 41022 34638 41074 34690
rect 42142 34638 42194 34690
rect 42814 34638 42866 34690
rect 43374 34638 43426 34690
rect 44382 34638 44434 34690
rect 49310 34638 49362 34690
rect 50654 34638 50706 34690
rect 51102 34638 51154 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 6526 34302 6578 34354
rect 11342 34302 11394 34354
rect 20526 34302 20578 34354
rect 24670 34302 24722 34354
rect 33406 34302 33458 34354
rect 33630 34302 33682 34354
rect 34302 34302 34354 34354
rect 35422 34302 35474 34354
rect 37886 34302 37938 34354
rect 38446 34302 38498 34354
rect 39566 34302 39618 34354
rect 50094 34302 50146 34354
rect 6750 34190 6802 34242
rect 7198 34190 7250 34242
rect 7422 34190 7474 34242
rect 7534 34190 7586 34242
rect 10110 34190 10162 34242
rect 13582 34190 13634 34242
rect 15598 34190 15650 34242
rect 19294 34190 19346 34242
rect 24334 34190 24386 34242
rect 33294 34190 33346 34242
rect 33966 34190 34018 34242
rect 34078 34190 34130 34242
rect 34862 34190 34914 34242
rect 38670 34190 38722 34242
rect 42926 34190 42978 34242
rect 44382 34190 44434 34242
rect 5294 34078 5346 34130
rect 6190 34078 6242 34130
rect 6414 34078 6466 34130
rect 6974 34078 7026 34130
rect 8990 34078 9042 34130
rect 12014 34078 12066 34130
rect 12574 34078 12626 34130
rect 12686 34078 12738 34130
rect 13022 34078 13074 34130
rect 15038 34078 15090 34130
rect 18622 34078 18674 34130
rect 19182 34078 19234 34130
rect 20862 34078 20914 34130
rect 27134 34078 27186 34130
rect 34526 34078 34578 34130
rect 38222 34078 38274 34130
rect 38558 34078 38610 34130
rect 38894 34078 38946 34130
rect 43038 34078 43090 34130
rect 43822 34078 43874 34130
rect 44158 34078 44210 34130
rect 49646 34078 49698 34130
rect 50318 34078 50370 34130
rect 50654 34078 50706 34130
rect 9998 33966 10050 34018
rect 10894 33966 10946 34018
rect 15598 33966 15650 34018
rect 21646 33966 21698 34018
rect 23774 33966 23826 34018
rect 27806 33966 27858 34018
rect 29934 33966 29986 34018
rect 30606 33966 30658 34018
rect 35758 33966 35810 34018
rect 42590 33966 42642 34018
rect 48862 33966 48914 34018
rect 50206 33966 50258 34018
rect 5518 33854 5570 33906
rect 5742 33854 5794 33906
rect 8878 33854 8930 33906
rect 9662 33854 9714 33906
rect 9774 33854 9826 33906
rect 53006 33854 53058 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 43486 33518 43538 33570
rect 50878 33518 50930 33570
rect 7982 33406 8034 33458
rect 9998 33406 10050 33458
rect 12910 33406 12962 33458
rect 16382 33406 16434 33458
rect 21982 33406 22034 33458
rect 24894 33406 24946 33458
rect 28254 33406 28306 33458
rect 29486 33406 29538 33458
rect 32846 33406 32898 33458
rect 33854 33406 33906 33458
rect 34414 33406 34466 33458
rect 44830 33406 44882 33458
rect 8318 33294 8370 33346
rect 9886 33294 9938 33346
rect 10222 33294 10274 33346
rect 11006 33294 11058 33346
rect 17390 33294 17442 33346
rect 21758 33294 21810 33346
rect 22094 33294 22146 33346
rect 22430 33294 22482 33346
rect 27806 33294 27858 33346
rect 31614 33294 31666 33346
rect 32398 33294 32450 33346
rect 41694 33294 41746 33346
rect 42142 33294 42194 33346
rect 42702 33294 42754 33346
rect 43150 33294 43202 33346
rect 45390 33294 45442 33346
rect 46062 33294 46114 33346
rect 48750 33294 48802 33346
rect 49422 33294 49474 33346
rect 27022 33182 27074 33234
rect 42030 33182 42082 33234
rect 49086 33182 49138 33234
rect 49758 33182 49810 33234
rect 8094 33070 8146 33122
rect 9214 33070 9266 33122
rect 11230 33070 11282 33122
rect 17950 33070 18002 33122
rect 37214 33070 37266 33122
rect 39902 33070 39954 33122
rect 45726 33070 45778 33122
rect 50206 33070 50258 33122
rect 50990 33070 51042 33122
rect 51102 33070 51154 33122
rect 51662 33070 51714 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 9662 32734 9714 32786
rect 21646 32734 21698 32786
rect 25566 32734 25618 32786
rect 26238 32734 26290 32786
rect 33518 32734 33570 32786
rect 36990 32734 37042 32786
rect 37550 32734 37602 32786
rect 38670 32734 38722 32786
rect 39118 32734 39170 32786
rect 39230 32734 39282 32786
rect 39902 32734 39954 32786
rect 42254 32734 42306 32786
rect 42590 32734 42642 32786
rect 43710 32734 43762 32786
rect 44494 32734 44546 32786
rect 45054 32734 45106 32786
rect 49310 32734 49362 32786
rect 49534 32734 49586 32786
rect 49870 32734 49922 32786
rect 50094 32734 50146 32786
rect 5742 32622 5794 32674
rect 14926 32622 14978 32674
rect 15150 32622 15202 32674
rect 15486 32622 15538 32674
rect 21870 32622 21922 32674
rect 25790 32622 25842 32674
rect 33406 32622 33458 32674
rect 42478 32622 42530 32674
rect 52446 32622 52498 32674
rect 1822 32510 1874 32562
rect 5630 32510 5682 32562
rect 5966 32510 6018 32562
rect 8766 32510 8818 32562
rect 15934 32510 15986 32562
rect 21982 32510 22034 32562
rect 25454 32510 25506 32562
rect 25902 32510 25954 32562
rect 26238 32510 26290 32562
rect 26574 32510 26626 32562
rect 33742 32510 33794 32562
rect 33966 32510 34018 32562
rect 37662 32510 37714 32562
rect 37774 32510 37826 32562
rect 37886 32510 37938 32562
rect 38110 32510 38162 32562
rect 38894 32510 38946 32562
rect 39342 32510 39394 32562
rect 39566 32510 39618 32562
rect 40126 32510 40178 32562
rect 41806 32510 41858 32562
rect 42030 32510 42082 32562
rect 43598 32510 43650 32562
rect 43934 32510 43986 32562
rect 44158 32510 44210 32562
rect 44942 32510 44994 32562
rect 45614 32510 45666 32562
rect 53118 32510 53170 32562
rect 2494 32398 2546 32450
rect 4622 32398 4674 32450
rect 5182 32398 5234 32450
rect 6414 32398 6466 32450
rect 15038 32398 15090 32450
rect 16270 32398 16322 32450
rect 27022 32398 27074 32450
rect 34750 32398 34802 32450
rect 43262 32398 43314 32450
rect 49086 32398 49138 32450
rect 49422 32398 49474 32450
rect 50318 32398 50370 32450
rect 45054 32286 45106 32338
rect 48862 32286 48914 32338
rect 49758 32286 49810 32338
rect 50094 32286 50146 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 15150 31950 15202 32002
rect 31726 31950 31778 32002
rect 37214 31950 37266 32002
rect 37550 31950 37602 32002
rect 50206 31950 50258 32002
rect 4958 31838 5010 31890
rect 5854 31838 5906 31890
rect 7870 31838 7922 31890
rect 9438 31838 9490 31890
rect 12686 31838 12738 31890
rect 13694 31838 13746 31890
rect 14478 31838 14530 31890
rect 25006 31838 25058 31890
rect 28478 31838 28530 31890
rect 31054 31838 31106 31890
rect 37662 31838 37714 31890
rect 38446 31838 38498 31890
rect 48526 31838 48578 31890
rect 50542 31838 50594 31890
rect 5070 31726 5122 31778
rect 5966 31726 6018 31778
rect 6302 31726 6354 31778
rect 7982 31726 8034 31778
rect 9774 31726 9826 31778
rect 13806 31726 13858 31778
rect 15038 31726 15090 31778
rect 16718 31726 16770 31778
rect 23662 31726 23714 31778
rect 24894 31726 24946 31778
rect 26350 31726 26402 31778
rect 26686 31726 26738 31778
rect 26910 31726 26962 31778
rect 27470 31726 27522 31778
rect 27918 31726 27970 31778
rect 28590 31726 28642 31778
rect 31390 31726 31442 31778
rect 32286 31726 32338 31778
rect 33966 31726 34018 31778
rect 34638 31726 34690 31778
rect 39006 31726 39058 31778
rect 39902 31726 39954 31778
rect 43374 31726 43426 31778
rect 45726 31726 45778 31778
rect 4734 31614 4786 31666
rect 5742 31614 5794 31666
rect 6862 31614 6914 31666
rect 10558 31614 10610 31666
rect 15598 31614 15650 31666
rect 16606 31614 16658 31666
rect 24670 31614 24722 31666
rect 27358 31614 27410 31666
rect 31614 31614 31666 31666
rect 31726 31614 31778 31666
rect 33406 31614 33458 31666
rect 40574 31614 40626 31666
rect 46398 31614 46450 31666
rect 6526 31502 6578 31554
rect 6750 31502 6802 31554
rect 7534 31502 7586 31554
rect 7758 31502 7810 31554
rect 23774 31502 23826 31554
rect 26014 31502 26066 31554
rect 26462 31502 26514 31554
rect 27246 31502 27298 31554
rect 28142 31502 28194 31554
rect 28366 31502 28418 31554
rect 29262 31502 29314 31554
rect 30830 31502 30882 31554
rect 31054 31502 31106 31554
rect 33070 31502 33122 31554
rect 34302 31502 34354 31554
rect 34526 31502 34578 31554
rect 37102 31502 37154 31554
rect 42814 31502 42866 31554
rect 48974 31502 49026 31554
rect 49870 31502 49922 31554
rect 50430 31502 50482 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 6638 31166 6690 31218
rect 7534 31166 7586 31218
rect 10110 31166 10162 31218
rect 17726 31166 17778 31218
rect 24334 31166 24386 31218
rect 26686 31166 26738 31218
rect 27358 31166 27410 31218
rect 30494 31166 30546 31218
rect 31054 31166 31106 31218
rect 31278 31166 31330 31218
rect 33966 31166 34018 31218
rect 34526 31166 34578 31218
rect 43822 31166 43874 31218
rect 44382 31166 44434 31218
rect 45278 31166 45330 31218
rect 6078 31054 6130 31106
rect 6190 31054 6242 31106
rect 20414 31054 20466 31106
rect 21646 31054 21698 31106
rect 22094 31054 22146 31106
rect 22542 31054 22594 31106
rect 22654 31054 22706 31106
rect 23438 31054 23490 31106
rect 24222 31054 24274 31106
rect 27582 31054 27634 31106
rect 31838 31054 31890 31106
rect 33630 31054 33682 31106
rect 33742 31054 33794 31106
rect 34302 31054 34354 31106
rect 35310 31054 35362 31106
rect 44830 31054 44882 31106
rect 45054 31054 45106 31106
rect 52446 31054 52498 31106
rect 6526 30942 6578 30994
rect 6750 30942 6802 30994
rect 7198 30942 7250 30994
rect 9774 30942 9826 30994
rect 9998 30942 10050 30994
rect 10222 30942 10274 30994
rect 16046 30942 16098 30994
rect 21086 30942 21138 30994
rect 21534 30942 21586 30994
rect 21758 30942 21810 30994
rect 22318 30942 22370 30994
rect 23550 30942 23602 30994
rect 24110 30942 24162 30994
rect 27694 30942 27746 30994
rect 28142 30942 28194 30994
rect 30830 30942 30882 30994
rect 31390 30942 31442 30994
rect 34190 30942 34242 30994
rect 45390 30942 45442 30994
rect 53118 30942 53170 30994
rect 13134 30830 13186 30882
rect 16382 30830 16434 30882
rect 16494 30830 16546 30882
rect 18286 30830 18338 30882
rect 34862 30830 34914 30882
rect 49982 30830 50034 30882
rect 50318 30830 50370 30882
rect 6078 30718 6130 30770
rect 7310 30718 7362 30770
rect 7534 30718 7586 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 9886 30382 9938 30434
rect 21982 30382 22034 30434
rect 31278 30382 31330 30434
rect 45166 30382 45218 30434
rect 4622 30270 4674 30322
rect 7198 30270 7250 30322
rect 15822 30270 15874 30322
rect 17950 30270 18002 30322
rect 24782 30270 24834 30322
rect 28590 30270 28642 30322
rect 43598 30270 43650 30322
rect 1710 30158 1762 30210
rect 5070 30158 5122 30210
rect 6414 30158 6466 30210
rect 9326 30158 9378 30210
rect 15486 30158 15538 30210
rect 16158 30158 16210 30210
rect 16942 30158 16994 30210
rect 18174 30158 18226 30210
rect 19406 30158 19458 30210
rect 22094 30158 22146 30210
rect 22318 30158 22370 30210
rect 22654 30158 22706 30210
rect 23886 30158 23938 30210
rect 25006 30158 25058 30210
rect 26126 30158 26178 30210
rect 29150 30158 29202 30210
rect 31390 30158 31442 30210
rect 42142 30158 42194 30210
rect 43150 30158 43202 30210
rect 43374 30158 43426 30210
rect 2494 30046 2546 30098
rect 6190 30046 6242 30098
rect 6302 30046 6354 30098
rect 6750 30046 6802 30098
rect 17278 30046 17330 30098
rect 18846 30046 18898 30098
rect 22542 30046 22594 30098
rect 23102 30046 23154 30098
rect 24558 30046 24610 30098
rect 25342 30046 25394 30098
rect 26462 30046 26514 30098
rect 29710 30046 29762 30098
rect 45278 30046 45330 30098
rect 52894 30046 52946 30098
rect 53230 30046 53282 30098
rect 9550 29934 9602 29986
rect 9774 29934 9826 29986
rect 21534 29934 21586 29986
rect 21982 29934 22034 29986
rect 23774 29934 23826 29986
rect 25678 29934 25730 29986
rect 26350 29934 26402 29986
rect 27022 29934 27074 29986
rect 28030 29934 28082 29986
rect 30270 29934 30322 29986
rect 31278 29934 31330 29986
rect 31950 29934 32002 29986
rect 39454 29934 39506 29986
rect 40574 29934 40626 29986
rect 42590 29934 42642 29986
rect 43598 29934 43650 29986
rect 43710 29934 43762 29986
rect 45166 29934 45218 29986
rect 45726 29934 45778 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 6862 29598 6914 29650
rect 9998 29598 10050 29650
rect 10110 29598 10162 29650
rect 12910 29598 12962 29650
rect 18958 29598 19010 29650
rect 26910 29598 26962 29650
rect 27918 29598 27970 29650
rect 31054 29598 31106 29650
rect 31502 29598 31554 29650
rect 31726 29598 31778 29650
rect 34190 29598 34242 29650
rect 35198 29598 35250 29650
rect 39230 29598 39282 29650
rect 41134 29598 41186 29650
rect 45502 29598 45554 29650
rect 53342 29598 53394 29650
rect 5854 29486 5906 29538
rect 8654 29486 8706 29538
rect 8878 29486 8930 29538
rect 9662 29486 9714 29538
rect 11902 29486 11954 29538
rect 18398 29486 18450 29538
rect 18846 29486 18898 29538
rect 20302 29486 20354 29538
rect 27806 29486 27858 29538
rect 30718 29486 30770 29538
rect 30830 29486 30882 29538
rect 31278 29486 31330 29538
rect 34526 29486 34578 29538
rect 34974 29486 35026 29538
rect 35534 29486 35586 29538
rect 40126 29486 40178 29538
rect 40350 29486 40402 29538
rect 47406 29486 47458 29538
rect 47854 29486 47906 29538
rect 48190 29486 48242 29538
rect 51214 29486 51266 29538
rect 6078 29374 6130 29426
rect 6414 29374 6466 29426
rect 6750 29374 6802 29426
rect 9886 29374 9938 29426
rect 10446 29374 10498 29426
rect 10782 29374 10834 29426
rect 11006 29374 11058 29426
rect 12126 29374 12178 29426
rect 13470 29374 13522 29426
rect 17726 29374 17778 29426
rect 18286 29374 18338 29426
rect 18734 29374 18786 29426
rect 20414 29374 20466 29426
rect 26798 29374 26850 29426
rect 28254 29374 28306 29426
rect 32174 29374 32226 29426
rect 34862 29374 34914 29426
rect 35982 29374 36034 29426
rect 39678 29374 39730 29426
rect 40798 29374 40850 29426
rect 41134 29374 41186 29426
rect 41358 29374 41410 29426
rect 42030 29374 42082 29426
rect 46510 29374 46562 29426
rect 46846 29374 46898 29426
rect 51886 29374 51938 29426
rect 52446 29374 52498 29426
rect 6190 29262 6242 29314
rect 8990 29262 9042 29314
rect 10894 29262 10946 29314
rect 12686 29262 12738 29314
rect 13022 29262 13074 29314
rect 14142 29262 14194 29314
rect 16270 29262 16322 29314
rect 16830 29262 16882 29314
rect 26462 29262 26514 29314
rect 28814 29262 28866 29314
rect 36654 29262 36706 29314
rect 38782 29262 38834 29314
rect 39902 29262 39954 29314
rect 42702 29262 42754 29314
rect 44830 29262 44882 29314
rect 49086 29262 49138 29314
rect 6638 29150 6690 29202
rect 31838 29150 31890 29202
rect 47070 29150 47122 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 6414 28814 6466 28866
rect 10110 28814 10162 28866
rect 11790 28814 11842 28866
rect 40798 28814 40850 28866
rect 47070 28814 47122 28866
rect 47406 28814 47458 28866
rect 10222 28702 10274 28754
rect 13694 28702 13746 28754
rect 16494 28702 16546 28754
rect 18286 28702 18338 28754
rect 18734 28702 18786 28754
rect 20302 28702 20354 28754
rect 20750 28702 20802 28754
rect 23214 28702 23266 28754
rect 27022 28702 27074 28754
rect 32174 28702 32226 28754
rect 34302 28702 34354 28754
rect 34974 28702 35026 28754
rect 35870 28702 35922 28754
rect 5742 28590 5794 28642
rect 8206 28590 8258 28642
rect 8430 28590 8482 28642
rect 8542 28590 8594 28642
rect 11454 28590 11506 28642
rect 12014 28590 12066 28642
rect 12910 28590 12962 28642
rect 17614 28590 17666 28642
rect 18174 28590 18226 28642
rect 19630 28590 19682 28642
rect 20078 28590 20130 28642
rect 27582 28590 27634 28642
rect 31390 28590 31442 28642
rect 36542 28590 36594 28642
rect 37214 28590 37266 28642
rect 37438 28590 37490 28642
rect 37550 28590 37602 28642
rect 37774 28590 37826 28642
rect 39678 28590 39730 28642
rect 40462 28590 40514 28642
rect 41358 28590 41410 28642
rect 47966 28590 48018 28642
rect 48190 28590 48242 28642
rect 48302 28590 48354 28642
rect 49086 28590 49138 28642
rect 49646 28590 49698 28642
rect 5854 28478 5906 28530
rect 5966 28478 6018 28530
rect 12798 28478 12850 28530
rect 22542 28478 22594 28530
rect 22654 28478 22706 28530
rect 30942 28478 30994 28530
rect 31054 28478 31106 28530
rect 36206 28478 36258 28530
rect 36318 28478 36370 28530
rect 36990 28478 37042 28530
rect 37998 28478 38050 28530
rect 38110 28478 38162 28530
rect 39342 28478 39394 28530
rect 40126 28478 40178 28530
rect 40686 28478 40738 28530
rect 41806 28478 41858 28530
rect 46510 28478 46562 28530
rect 46734 28478 46786 28530
rect 8990 28366 9042 28418
rect 22878 28366 22930 28418
rect 28030 28366 28082 28418
rect 30494 28366 30546 28418
rect 30718 28366 30770 28418
rect 39006 28366 39058 28418
rect 39454 28366 39506 28418
rect 40238 28366 40290 28418
rect 40798 28366 40850 28418
rect 48750 28366 48802 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 5294 27918 5346 27970
rect 5966 27974 6018 28026
rect 6190 28030 6242 28082
rect 7534 28030 7586 28082
rect 8318 28030 8370 28082
rect 21758 28030 21810 28082
rect 22766 28030 22818 28082
rect 23886 28030 23938 28082
rect 24670 28030 24722 28082
rect 34190 28030 34242 28082
rect 34526 28030 34578 28082
rect 34974 28030 35026 28082
rect 35534 28030 35586 28082
rect 35982 28030 36034 28082
rect 36766 28030 36818 28082
rect 40238 28030 40290 28082
rect 40462 28030 40514 28082
rect 41022 28030 41074 28082
rect 45390 28030 45442 28082
rect 46734 28030 46786 28082
rect 47630 28030 47682 28082
rect 48078 28030 48130 28082
rect 48974 28030 49026 28082
rect 6638 27918 6690 27970
rect 7310 27918 7362 27970
rect 7758 27918 7810 27970
rect 10334 27918 10386 27970
rect 10670 27918 10722 27970
rect 19742 27918 19794 27970
rect 21870 27918 21922 27970
rect 23102 27918 23154 27970
rect 23438 27918 23490 27970
rect 24110 27918 24162 27970
rect 31278 27918 31330 27970
rect 34862 27918 34914 27970
rect 45614 27918 45666 27970
rect 46510 27918 46562 27970
rect 1710 27806 1762 27858
rect 4958 27806 5010 27858
rect 5854 27806 5906 27858
rect 6526 27806 6578 27858
rect 6974 27806 7026 27858
rect 7198 27806 7250 27858
rect 19070 27806 19122 27858
rect 19630 27806 19682 27858
rect 20190 27806 20242 27858
rect 21534 27806 21586 27858
rect 23550 27806 23602 27858
rect 24222 27806 24274 27858
rect 27246 27806 27298 27858
rect 40126 27806 40178 27858
rect 44270 27806 44322 27858
rect 45054 27806 45106 27858
rect 45726 27806 45778 27858
rect 46398 27806 46450 27858
rect 53118 27806 53170 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 6862 27694 6914 27746
rect 23214 27694 23266 27746
rect 26910 27694 26962 27746
rect 44606 27694 44658 27746
rect 49982 27694 50034 27746
rect 50318 27694 50370 27746
rect 52446 27694 52498 27746
rect 34974 27582 35026 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 6638 27246 6690 27298
rect 27582 27246 27634 27298
rect 37102 27246 37154 27298
rect 45054 27246 45106 27298
rect 45390 27246 45442 27298
rect 45726 27246 45778 27298
rect 46398 27246 46450 27298
rect 47518 27246 47570 27298
rect 4846 27134 4898 27186
rect 6526 27134 6578 27186
rect 16382 27134 16434 27186
rect 16830 27134 16882 27186
rect 23886 27134 23938 27186
rect 26014 27134 26066 27186
rect 32286 27134 32338 27186
rect 32734 27134 32786 27186
rect 45950 27134 46002 27186
rect 47630 27134 47682 27186
rect 11006 27022 11058 27074
rect 11342 27022 11394 27074
rect 11678 27022 11730 27074
rect 12238 27022 12290 27074
rect 12462 27022 12514 27074
rect 13470 27022 13522 27074
rect 21422 27022 21474 27074
rect 21646 27022 21698 27074
rect 21982 27022 22034 27074
rect 23102 27022 23154 27074
rect 30494 27022 30546 27074
rect 31278 27022 31330 27074
rect 31838 27022 31890 27074
rect 34526 27022 34578 27074
rect 35086 27022 35138 27074
rect 35646 27022 35698 27074
rect 36318 27022 36370 27074
rect 37214 27022 37266 27074
rect 38446 27022 38498 27074
rect 39118 27022 39170 27074
rect 40238 27022 40290 27074
rect 40686 27022 40738 27074
rect 41470 27022 41522 27074
rect 44830 27022 44882 27074
rect 46622 27022 46674 27074
rect 47070 27022 47122 27074
rect 53230 27022 53282 27074
rect 14254 26910 14306 26962
rect 22206 26910 22258 26962
rect 22542 26910 22594 26962
rect 27694 26910 27746 26962
rect 30606 26910 30658 26962
rect 30718 26910 30770 26962
rect 30830 26910 30882 26962
rect 31726 26910 31778 26962
rect 34862 26910 34914 26962
rect 35870 26910 35922 26962
rect 37662 26910 37714 26962
rect 37998 26910 38050 26962
rect 38670 26910 38722 26962
rect 39342 26910 39394 26962
rect 40014 26910 40066 26962
rect 41022 26910 41074 26962
rect 44270 26910 44322 26962
rect 52894 26910 52946 26962
rect 11230 26798 11282 26850
rect 11902 26798 11954 26850
rect 12014 26798 12066 26850
rect 21534 26798 21586 26850
rect 22430 26798 22482 26850
rect 27582 26798 27634 26850
rect 28142 26798 28194 26850
rect 31502 26798 31554 26850
rect 37102 26798 37154 26850
rect 37886 26798 37938 26850
rect 40126 26798 40178 26850
rect 48078 26798 48130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 6638 26462 6690 26514
rect 9550 26462 9602 26514
rect 11678 26462 11730 26514
rect 15598 26462 15650 26514
rect 24110 26462 24162 26514
rect 26798 26462 26850 26514
rect 30942 26462 30994 26514
rect 49198 26462 49250 26514
rect 51662 26462 51714 26514
rect 53342 26462 53394 26514
rect 5742 26350 5794 26402
rect 6078 26350 6130 26402
rect 12910 26350 12962 26402
rect 15262 26350 15314 26402
rect 29038 26350 29090 26402
rect 31166 26350 31218 26402
rect 45166 26350 45218 26402
rect 49870 26350 49922 26402
rect 6526 26238 6578 26290
rect 6750 26238 6802 26290
rect 7198 26238 7250 26290
rect 9774 26238 9826 26290
rect 11342 26238 11394 26290
rect 11566 26238 11618 26290
rect 11790 26238 11842 26290
rect 11902 26238 11954 26290
rect 12350 26238 12402 26290
rect 12574 26238 12626 26290
rect 17726 26238 17778 26290
rect 18286 26238 18338 26290
rect 24446 26238 24498 26290
rect 29822 26238 29874 26290
rect 31390 26238 31442 26290
rect 31614 26238 31666 26290
rect 37774 26238 37826 26290
rect 39678 26238 39730 26290
rect 40126 26238 40178 26290
rect 40238 26238 40290 26290
rect 43822 26238 43874 26290
rect 44606 26238 44658 26290
rect 49086 26238 49138 26290
rect 49758 26238 49810 26290
rect 51214 26238 51266 26290
rect 51886 26238 51938 26290
rect 13358 26126 13410 26178
rect 18398 26126 18450 26178
rect 18846 26126 18898 26178
rect 22766 26126 22818 26178
rect 30270 26126 30322 26178
rect 31726 26126 31778 26178
rect 32174 26126 32226 26178
rect 39902 26126 39954 26178
rect 40910 26126 40962 26178
rect 43038 26126 43090 26178
rect 44270 26126 44322 26178
rect 12798 26014 12850 26066
rect 13134 26014 13186 26066
rect 13358 26014 13410 26066
rect 37998 26014 38050 26066
rect 38334 26014 38386 26066
rect 49198 26014 49250 26066
rect 49870 26014 49922 26066
rect 51550 26014 51602 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6974 25678 7026 25730
rect 19294 25678 19346 25730
rect 19630 25678 19682 25730
rect 34862 25678 34914 25730
rect 35198 25678 35250 25730
rect 6638 25566 6690 25618
rect 31950 25566 32002 25618
rect 34190 25566 34242 25618
rect 35198 25566 35250 25618
rect 5630 25454 5682 25506
rect 5854 25454 5906 25506
rect 6078 25454 6130 25506
rect 6302 25454 6354 25506
rect 8990 25454 9042 25506
rect 17950 25454 18002 25506
rect 18398 25454 18450 25506
rect 18622 25454 18674 25506
rect 19070 25454 19122 25506
rect 19518 25454 19570 25506
rect 25902 25454 25954 25506
rect 26574 25454 26626 25506
rect 27694 25454 27746 25506
rect 27918 25454 27970 25506
rect 28142 25454 28194 25506
rect 29374 25454 29426 25506
rect 31278 25454 31330 25506
rect 49198 25454 49250 25506
rect 49870 25454 49922 25506
rect 50878 25454 50930 25506
rect 51102 25454 51154 25506
rect 51662 25454 51714 25506
rect 6750 25342 6802 25394
rect 9438 25342 9490 25394
rect 9662 25342 9714 25394
rect 10334 25342 10386 25394
rect 10670 25342 10722 25394
rect 18958 25342 19010 25394
rect 26238 25342 26290 25394
rect 26910 25342 26962 25394
rect 29150 25342 29202 25394
rect 29934 25342 29986 25394
rect 49646 25342 49698 25394
rect 50206 25342 50258 25394
rect 50430 25342 50482 25394
rect 51326 25342 51378 25394
rect 53230 25342 53282 25394
rect 5966 25230 6018 25282
rect 8990 25230 9042 25282
rect 25566 25230 25618 25282
rect 26798 25230 26850 25282
rect 28478 25230 28530 25282
rect 30382 25230 30434 25282
rect 34750 25230 34802 25282
rect 43374 25230 43426 25282
rect 48414 25230 48466 25282
rect 49534 25230 49586 25282
rect 50542 25230 50594 25282
rect 51550 25230 51602 25282
rect 52894 25230 52946 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 5070 24894 5122 24946
rect 5966 24894 6018 24946
rect 6974 24894 7026 24946
rect 11454 24894 11506 24946
rect 13134 24894 13186 24946
rect 18510 24894 18562 24946
rect 19070 24894 19122 24946
rect 29150 24894 29202 24946
rect 30270 24894 30322 24946
rect 34974 24894 35026 24946
rect 42478 24894 42530 24946
rect 43710 24894 43762 24946
rect 49086 24894 49138 24946
rect 50654 24894 50706 24946
rect 51550 24894 51602 24946
rect 11678 24782 11730 24834
rect 12350 24782 12402 24834
rect 13582 24782 13634 24834
rect 18622 24782 18674 24834
rect 22318 24782 22370 24834
rect 26126 24782 26178 24834
rect 28366 24782 28418 24834
rect 28590 24782 28642 24834
rect 29710 24782 29762 24834
rect 34414 24782 34466 24834
rect 34750 24782 34802 24834
rect 48862 24782 48914 24834
rect 50878 24782 50930 24834
rect 1710 24670 1762 24722
rect 5406 24670 5458 24722
rect 5630 24670 5682 24722
rect 6638 24670 6690 24722
rect 11342 24670 11394 24722
rect 11790 24670 11842 24722
rect 12686 24670 12738 24722
rect 13134 24670 13186 24722
rect 13470 24670 13522 24722
rect 18286 24670 18338 24722
rect 22990 24670 23042 24722
rect 26462 24670 26514 24722
rect 26910 24670 26962 24722
rect 29038 24670 29090 24722
rect 29598 24670 29650 24722
rect 30718 24670 30770 24722
rect 34526 24670 34578 24722
rect 35534 24670 35586 24722
rect 39006 24670 39058 24722
rect 40350 24670 40402 24722
rect 42702 24670 42754 24722
rect 42926 24670 42978 24722
rect 45390 24670 45442 24722
rect 48750 24670 48802 24722
rect 49422 24670 49474 24722
rect 50542 24670 50594 24722
rect 51438 24670 51490 24722
rect 51662 24670 51714 24722
rect 51886 24670 51938 24722
rect 53230 24670 53282 24722
rect 2494 24558 2546 24610
rect 4622 24558 4674 24610
rect 11678 24558 11730 24610
rect 12798 24558 12850 24610
rect 20078 24558 20130 24610
rect 23662 24558 23714 24610
rect 26238 24558 26290 24610
rect 27470 24558 27522 24610
rect 28142 24558 28194 24610
rect 34638 24558 34690 24610
rect 36206 24558 36258 24610
rect 38334 24558 38386 24610
rect 39342 24558 39394 24610
rect 39790 24558 39842 24610
rect 42366 24558 42418 24610
rect 44270 24558 44322 24610
rect 44830 24558 44882 24610
rect 46062 24558 46114 24610
rect 48190 24558 48242 24610
rect 50206 24558 50258 24610
rect 26686 24446 26738 24498
rect 28926 24446 28978 24498
rect 29486 24446 29538 24498
rect 44046 24446 44098 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 2606 24110 2658 24162
rect 2942 24110 2994 24162
rect 46622 24110 46674 24162
rect 46958 24110 47010 24162
rect 14702 23998 14754 24050
rect 16830 23998 16882 24050
rect 17278 23998 17330 24050
rect 19070 23998 19122 24050
rect 22542 23998 22594 24050
rect 24782 23998 24834 24050
rect 27134 23998 27186 24050
rect 29934 23998 29986 24050
rect 32062 23998 32114 24050
rect 36206 23998 36258 24050
rect 38782 23998 38834 24050
rect 40798 23998 40850 24050
rect 43822 23998 43874 24050
rect 44942 23998 44994 24050
rect 49870 23998 49922 24050
rect 7870 23886 7922 23938
rect 11790 23886 11842 23938
rect 13918 23886 13970 23938
rect 18510 23886 18562 23938
rect 18958 23886 19010 23938
rect 25566 23886 25618 23938
rect 29262 23886 29314 23938
rect 34638 23886 34690 23938
rect 34974 23886 35026 23938
rect 35646 23886 35698 23938
rect 36318 23886 36370 23938
rect 37214 23886 37266 23938
rect 41358 23886 41410 23938
rect 43038 23886 43090 23938
rect 44270 23886 44322 23938
rect 45278 23886 45330 23938
rect 50430 23886 50482 23938
rect 5630 23774 5682 23826
rect 11566 23774 11618 23826
rect 35982 23774 36034 23826
rect 36094 23774 36146 23826
rect 36878 23774 36930 23826
rect 42142 23774 42194 23826
rect 46286 23774 46338 23826
rect 46734 23774 46786 23826
rect 50318 23774 50370 23826
rect 2718 23662 2770 23714
rect 3502 23662 3554 23714
rect 5966 23662 6018 23714
rect 8094 23662 8146 23714
rect 26014 23662 26066 23714
rect 28590 23662 28642 23714
rect 34862 23662 34914 23714
rect 37102 23662 37154 23714
rect 45614 23662 45666 23714
rect 48190 23662 48242 23714
rect 50094 23662 50146 23714
rect 50878 23662 50930 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 6414 23326 6466 23378
rect 11230 23326 11282 23378
rect 11454 23326 11506 23378
rect 31614 23326 31666 23378
rect 36542 23326 36594 23378
rect 37214 23326 37266 23378
rect 37774 23326 37826 23378
rect 41246 23326 41298 23378
rect 43598 23326 43650 23378
rect 49310 23326 49362 23378
rect 49758 23326 49810 23378
rect 4846 23214 4898 23266
rect 5070 23214 5122 23266
rect 10110 23214 10162 23266
rect 12686 23214 12738 23266
rect 20078 23214 20130 23266
rect 20414 23214 20466 23266
rect 39454 23214 39506 23266
rect 6190 23102 6242 23154
rect 10446 23102 10498 23154
rect 10670 23102 10722 23154
rect 10894 23102 10946 23154
rect 13022 23102 13074 23154
rect 19518 23102 19570 23154
rect 20638 23102 20690 23154
rect 21198 23102 21250 23154
rect 31502 23102 31554 23154
rect 37102 23102 37154 23154
rect 41246 23102 41298 23154
rect 41582 23102 41634 23154
rect 42030 23102 42082 23154
rect 43934 23102 43986 23154
rect 44046 23102 44098 23154
rect 44942 23102 44994 23154
rect 48750 23102 48802 23154
rect 49646 23102 49698 23154
rect 53118 23102 53170 23154
rect 4622 22990 4674 23042
rect 10558 22990 10610 23042
rect 27358 22990 27410 23042
rect 39342 22990 39394 23042
rect 42590 22990 42642 23042
rect 43486 22990 43538 23042
rect 45390 22990 45442 23042
rect 47966 22990 48018 23042
rect 50318 22990 50370 23042
rect 52446 22990 52498 23042
rect 5182 22878 5234 22930
rect 11566 22878 11618 22930
rect 13022 22878 13074 22930
rect 37214 22878 37266 22930
rect 39678 22878 39730 22930
rect 49758 22878 49810 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 8318 22542 8370 22594
rect 8990 22542 9042 22594
rect 9550 22542 9602 22594
rect 10558 22542 10610 22594
rect 15934 22542 15986 22594
rect 4622 22430 4674 22482
rect 5070 22430 5122 22482
rect 7086 22430 7138 22482
rect 9326 22430 9378 22482
rect 13694 22430 13746 22482
rect 18286 22430 18338 22482
rect 27134 22430 27186 22482
rect 29934 22430 29986 22482
rect 31502 22430 31554 22482
rect 32622 22430 32674 22482
rect 34750 22430 34802 22482
rect 41806 22430 41858 22482
rect 43038 22430 43090 22482
rect 47742 22430 47794 22482
rect 49198 22430 49250 22482
rect 52782 22430 52834 22482
rect 1710 22318 1762 22370
rect 8318 22318 8370 22370
rect 8766 22318 8818 22370
rect 9438 22318 9490 22370
rect 10222 22318 10274 22370
rect 10782 22318 10834 22370
rect 13918 22318 13970 22370
rect 14030 22318 14082 22370
rect 14366 22318 14418 22370
rect 14814 22318 14866 22370
rect 24334 22318 24386 22370
rect 27358 22318 27410 22370
rect 27694 22318 27746 22370
rect 28030 22318 28082 22370
rect 29486 22318 29538 22370
rect 31838 22318 31890 22370
rect 37998 22318 38050 22370
rect 39118 22318 39170 22370
rect 41134 22318 41186 22370
rect 42478 22318 42530 22370
rect 44830 22318 44882 22370
rect 48078 22318 48130 22370
rect 51326 22318 51378 22370
rect 2494 22206 2546 22258
rect 5854 22206 5906 22258
rect 6302 22206 6354 22258
rect 7422 22206 7474 22258
rect 7534 22206 7586 22258
rect 7758 22206 7810 22258
rect 7982 22206 8034 22258
rect 9998 22206 10050 22258
rect 13470 22206 13522 22258
rect 16046 22206 16098 22258
rect 18958 22206 19010 22258
rect 25006 22206 25058 22258
rect 27582 22206 27634 22258
rect 37326 22206 37378 22258
rect 40574 22206 40626 22258
rect 42142 22206 42194 22258
rect 45614 22206 45666 22258
rect 50990 22206 51042 22258
rect 51438 22206 51490 22258
rect 51550 22206 51602 22258
rect 52670 22206 52722 22258
rect 5742 22094 5794 22146
rect 5966 22094 6018 22146
rect 6078 22094 6130 22146
rect 10782 22094 10834 22146
rect 14030 22094 14082 22146
rect 17726 22094 17778 22146
rect 18622 22094 18674 22146
rect 30382 22094 30434 22146
rect 36430 22094 36482 22146
rect 41582 22094 41634 22146
rect 43598 22094 43650 22146
rect 44046 22094 44098 22146
rect 52110 22094 52162 22146
rect 52894 22094 52946 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 5406 21758 5458 21810
rect 5742 21758 5794 21810
rect 9550 21758 9602 21810
rect 16830 21758 16882 21810
rect 23886 21758 23938 21810
rect 26910 21758 26962 21810
rect 27134 21758 27186 21810
rect 27582 21758 27634 21810
rect 49982 21758 50034 21810
rect 2718 21646 2770 21698
rect 2942 21646 2994 21698
rect 5854 21646 5906 21698
rect 7310 21646 7362 21698
rect 7422 21646 7474 21698
rect 9662 21646 9714 21698
rect 14254 21646 14306 21698
rect 35310 21646 35362 21698
rect 39790 21646 39842 21698
rect 42366 21646 42418 21698
rect 50430 21646 50482 21698
rect 52670 21646 52722 21698
rect 52894 21646 52946 21698
rect 53230 21646 53282 21698
rect 5630 21534 5682 21586
rect 6526 21534 6578 21586
rect 6638 21534 6690 21586
rect 7086 21534 7138 21586
rect 13582 21534 13634 21586
rect 17726 21534 17778 21586
rect 20638 21534 20690 21586
rect 23998 21534 24050 21586
rect 24334 21534 24386 21586
rect 26798 21534 26850 21586
rect 34862 21534 34914 21586
rect 37102 21534 37154 21586
rect 37774 21534 37826 21586
rect 38110 21534 38162 21586
rect 38670 21534 38722 21586
rect 40238 21534 40290 21586
rect 41582 21534 41634 21586
rect 41806 21534 41858 21586
rect 42814 21534 42866 21586
rect 43150 21534 43202 21586
rect 44046 21534 44098 21586
rect 44494 21534 44546 21586
rect 49758 21534 49810 21586
rect 2606 21422 2658 21474
rect 3390 21422 3442 21474
rect 4846 21422 4898 21474
rect 6302 21422 6354 21474
rect 16382 21422 16434 21474
rect 18286 21422 18338 21474
rect 21310 21422 21362 21474
rect 23438 21422 23490 21474
rect 6190 21310 6242 21362
rect 23886 21310 23938 21362
rect 50094 21534 50146 21586
rect 24446 21422 24498 21474
rect 30718 21422 30770 21474
rect 34302 21422 34354 21474
rect 36206 21422 36258 21474
rect 41246 21422 41298 21474
rect 42702 21422 42754 21474
rect 45054 21422 45106 21474
rect 47742 21422 47794 21474
rect 24446 21310 24498 21362
rect 41022 21310 41074 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 6638 20974 6690 21026
rect 43710 20974 43762 21026
rect 43934 20974 43986 21026
rect 6526 20862 6578 20914
rect 10782 20862 10834 20914
rect 12910 20862 12962 20914
rect 29934 20862 29986 20914
rect 32958 20862 33010 20914
rect 42030 20862 42082 20914
rect 43598 20862 43650 20914
rect 5630 20750 5682 20802
rect 6190 20750 6242 20802
rect 9998 20750 10050 20802
rect 16830 20750 16882 20802
rect 23886 20750 23938 20802
rect 30382 20750 30434 20802
rect 31166 20750 31218 20802
rect 31838 20750 31890 20802
rect 33518 20750 33570 20802
rect 34862 20750 34914 20802
rect 37998 20750 38050 20802
rect 39118 20750 39170 20802
rect 41470 20750 41522 20802
rect 42142 20750 42194 20802
rect 42478 20750 42530 20802
rect 44942 20750 44994 20802
rect 45166 20750 45218 20802
rect 45390 20750 45442 20802
rect 45950 20750 46002 20802
rect 5966 20638 6018 20690
rect 23214 20638 23266 20690
rect 23438 20638 23490 20690
rect 29150 20638 29202 20690
rect 30830 20638 30882 20690
rect 32062 20638 32114 20690
rect 37326 20638 37378 20690
rect 40574 20638 40626 20690
rect 5742 20526 5794 20578
rect 9662 20526 9714 20578
rect 16606 20526 16658 20578
rect 23550 20526 23602 20578
rect 29262 20526 29314 20578
rect 29486 20526 29538 20578
rect 30942 20526 30994 20578
rect 31502 20526 31554 20578
rect 34526 20526 34578 20578
rect 41582 20526 41634 20578
rect 41694 20526 41746 20578
rect 43934 20526 43986 20578
rect 45054 20526 45106 20578
rect 49534 20526 49586 20578
rect 49870 20526 49922 20578
rect 50430 20526 50482 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 5854 20190 5906 20242
rect 41918 20190 41970 20242
rect 42254 20190 42306 20242
rect 47406 20190 47458 20242
rect 2830 20078 2882 20130
rect 3054 20078 3106 20130
rect 3502 20078 3554 20130
rect 7870 20078 7922 20130
rect 8094 20078 8146 20130
rect 9550 20078 9602 20130
rect 14702 20078 14754 20130
rect 15038 20078 15090 20130
rect 15374 20078 15426 20130
rect 15710 20078 15762 20130
rect 16494 20078 16546 20130
rect 16830 20078 16882 20130
rect 23998 20078 24050 20130
rect 26798 20078 26850 20130
rect 30494 20078 30546 20130
rect 31838 20078 31890 20130
rect 33182 20078 33234 20130
rect 37214 20078 37266 20130
rect 37438 20078 37490 20130
rect 40126 20078 40178 20130
rect 41806 20078 41858 20130
rect 42814 20078 42866 20130
rect 44046 20078 44098 20130
rect 44606 20078 44658 20130
rect 44830 20078 44882 20130
rect 45390 20078 45442 20130
rect 45502 20078 45554 20130
rect 46734 20078 46786 20130
rect 46958 20078 47010 20130
rect 47518 20078 47570 20130
rect 48862 20078 48914 20130
rect 49758 20078 49810 20130
rect 5182 19966 5234 20018
rect 5630 19966 5682 20018
rect 8206 19966 8258 20018
rect 9886 19966 9938 20018
rect 10334 19966 10386 20018
rect 10558 19966 10610 20018
rect 17502 19966 17554 20018
rect 20750 19966 20802 20018
rect 23774 19966 23826 20018
rect 24110 19966 24162 20018
rect 26126 19966 26178 20018
rect 26574 19966 26626 20018
rect 30270 19966 30322 20018
rect 32174 19966 32226 20018
rect 32398 19966 32450 20018
rect 37102 19966 37154 20018
rect 39790 19966 39842 20018
rect 40014 19966 40066 20018
rect 41470 19966 41522 20018
rect 43822 19966 43874 20018
rect 44494 19966 44546 20018
rect 44942 19966 44994 20018
rect 45614 19966 45666 20018
rect 46286 19966 46338 20018
rect 47294 19966 47346 20018
rect 48078 19966 48130 20018
rect 49422 19966 49474 20018
rect 50318 19966 50370 20018
rect 8654 19854 8706 19906
rect 11118 19854 11170 19906
rect 16270 19854 16322 19906
rect 18174 19854 18226 19906
rect 20302 19854 20354 19906
rect 21422 19854 21474 19906
rect 23550 19854 23602 19906
rect 24558 19854 24610 19906
rect 30942 19854 30994 19906
rect 33070 19854 33122 19906
rect 37886 19854 37938 19906
rect 41022 19854 41074 19906
rect 42366 19854 42418 19906
rect 43486 19854 43538 19906
rect 46062 19854 46114 19906
rect 46510 19854 46562 19906
rect 51102 19854 51154 19906
rect 53230 19854 53282 19906
rect 2718 19742 2770 19794
rect 10222 19742 10274 19794
rect 33406 19742 33458 19794
rect 37550 19742 37602 19794
rect 37886 19742 37938 19794
rect 47854 19742 47906 19794
rect 48750 19742 48802 19794
rect 49086 19742 49138 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 8430 19406 8482 19458
rect 8766 19406 8818 19458
rect 2494 19294 2546 19346
rect 4622 19294 4674 19346
rect 5182 19294 5234 19346
rect 11678 19294 11730 19346
rect 17054 19294 17106 19346
rect 23886 19294 23938 19346
rect 32846 19294 32898 19346
rect 37214 19294 37266 19346
rect 39230 19294 39282 19346
rect 47070 19294 47122 19346
rect 49310 19294 49362 19346
rect 52222 19294 52274 19346
rect 1710 19182 1762 19234
rect 11790 19182 11842 19234
rect 20526 19182 20578 19234
rect 23326 19182 23378 19234
rect 23774 19182 23826 19234
rect 23998 19182 24050 19234
rect 25454 19182 25506 19234
rect 29374 19182 29426 19234
rect 30270 19182 30322 19234
rect 33630 19182 33682 19234
rect 37550 19182 37602 19234
rect 41246 19182 41298 19234
rect 41582 19182 41634 19234
rect 48190 19182 48242 19234
rect 53230 19182 53282 19234
rect 11454 19070 11506 19122
rect 24334 19070 24386 19122
rect 26238 19070 26290 19122
rect 37998 19070 38050 19122
rect 39566 19070 39618 19122
rect 42142 19070 42194 19122
rect 47742 19070 47794 19122
rect 8654 18958 8706 19010
rect 20190 18958 20242 19010
rect 23102 18958 23154 19010
rect 24782 18958 24834 19010
rect 25118 18958 25170 19010
rect 28478 18958 28530 19010
rect 29038 18958 29090 19010
rect 29262 18958 29314 19010
rect 29822 18958 29874 19010
rect 33742 18958 33794 19010
rect 33966 18958 34018 19010
rect 34302 18958 34354 19010
rect 38782 18958 38834 19010
rect 40574 18958 40626 19010
rect 43822 18958 43874 19010
rect 44270 18958 44322 19010
rect 44942 18958 44994 19010
rect 45390 18958 45442 19010
rect 47406 18958 47458 19010
rect 52894 18958 52946 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 24558 18622 24610 18674
rect 32398 18622 32450 18674
rect 50990 18622 51042 18674
rect 6078 18510 6130 18562
rect 7982 18510 8034 18562
rect 8766 18510 8818 18562
rect 27134 18510 27186 18562
rect 31390 18510 31442 18562
rect 31726 18510 31778 18562
rect 31950 18510 32002 18562
rect 32510 18510 32562 18562
rect 38110 18510 38162 18562
rect 39118 18510 39170 18562
rect 40126 18510 40178 18562
rect 41246 18510 41298 18562
rect 43822 18510 43874 18562
rect 46622 18510 46674 18562
rect 49646 18510 49698 18562
rect 51438 18510 51490 18562
rect 6750 18398 6802 18450
rect 7534 18398 7586 18450
rect 8318 18398 8370 18450
rect 8990 18398 9042 18450
rect 12574 18398 12626 18450
rect 16270 18398 16322 18450
rect 26910 18398 26962 18450
rect 27022 18398 27074 18450
rect 27582 18398 27634 18450
rect 31502 18398 31554 18450
rect 32174 18398 32226 18450
rect 33182 18398 33234 18450
rect 37102 18398 37154 18450
rect 38446 18398 38498 18450
rect 38894 18398 38946 18450
rect 39790 18398 39842 18450
rect 41470 18398 41522 18450
rect 41694 18398 41746 18450
rect 41918 18398 41970 18450
rect 42590 18398 42642 18450
rect 43150 18398 43202 18450
rect 43486 18398 43538 18450
rect 45166 18398 45218 18450
rect 46958 18398 47010 18450
rect 49422 18398 49474 18450
rect 50766 18398 50818 18450
rect 51774 18398 51826 18450
rect 51886 18398 51938 18450
rect 52222 18398 52274 18450
rect 52446 18398 52498 18450
rect 52558 18398 52610 18450
rect 52894 18398 52946 18450
rect 6638 18286 6690 18338
rect 8654 18286 8706 18338
rect 9662 18286 9714 18338
rect 13246 18286 13298 18338
rect 15374 18286 15426 18338
rect 15710 18286 15762 18338
rect 25342 18286 25394 18338
rect 26574 18286 26626 18338
rect 31614 18286 31666 18338
rect 33854 18286 33906 18338
rect 35982 18286 36034 18338
rect 37438 18286 37490 18338
rect 37774 18286 37826 18338
rect 40238 18286 40290 18338
rect 44606 18286 44658 18338
rect 46734 18286 46786 18338
rect 47854 18286 47906 18338
rect 51550 18286 51602 18338
rect 15822 18174 15874 18226
rect 38446 18174 38498 18226
rect 42366 18174 42418 18226
rect 51102 18174 51154 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 9886 17838 9938 17890
rect 32622 17838 32674 17890
rect 42478 17838 42530 17890
rect 51214 17838 51266 17890
rect 9102 17726 9154 17778
rect 10110 17726 10162 17778
rect 10670 17726 10722 17778
rect 20750 17726 20802 17778
rect 29934 17726 29986 17778
rect 33630 17726 33682 17778
rect 36542 17726 36594 17778
rect 40686 17726 40738 17778
rect 43710 17726 43762 17778
rect 46622 17726 46674 17778
rect 48750 17726 48802 17778
rect 5630 17614 5682 17666
rect 5854 17614 5906 17666
rect 6190 17614 6242 17666
rect 6862 17614 6914 17666
rect 7422 17614 7474 17666
rect 8654 17614 8706 17666
rect 9662 17614 9714 17666
rect 17838 17614 17890 17666
rect 29150 17614 29202 17666
rect 33966 17614 34018 17666
rect 34414 17614 34466 17666
rect 39006 17614 39058 17666
rect 39566 17614 39618 17666
rect 43150 17614 43202 17666
rect 45950 17614 46002 17666
rect 49198 17614 49250 17666
rect 51998 17614 52050 17666
rect 6526 17502 6578 17554
rect 10222 17502 10274 17554
rect 18622 17502 18674 17554
rect 25790 17502 25842 17554
rect 32734 17502 32786 17554
rect 33182 17502 33234 17554
rect 33854 17502 33906 17554
rect 39230 17502 39282 17554
rect 42590 17502 42642 17554
rect 44158 17502 44210 17554
rect 50542 17502 50594 17554
rect 50654 17502 50706 17554
rect 51102 17502 51154 17554
rect 51214 17502 51266 17554
rect 51662 17502 51714 17554
rect 51774 17502 51826 17554
rect 6638 17390 6690 17442
rect 7086 17390 7138 17442
rect 8318 17390 8370 17442
rect 17054 17390 17106 17442
rect 17502 17390 17554 17442
rect 24894 17390 24946 17442
rect 25454 17390 25506 17442
rect 25678 17390 25730 17442
rect 28590 17390 28642 17442
rect 32174 17390 32226 17442
rect 34190 17390 34242 17442
rect 38110 17390 38162 17442
rect 38558 17390 38610 17442
rect 42926 17390 42978 17442
rect 44942 17390 44994 17442
rect 45502 17390 45554 17442
rect 50878 17390 50930 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 6414 17054 6466 17106
rect 7534 17054 7586 17106
rect 13134 17054 13186 17106
rect 15822 17054 15874 17106
rect 18174 17054 18226 17106
rect 24222 17054 24274 17106
rect 32286 17054 32338 17106
rect 36430 17054 36482 17106
rect 37998 17054 38050 17106
rect 51326 17054 51378 17106
rect 51774 17054 51826 17106
rect 2494 16942 2546 16994
rect 13918 16942 13970 16994
rect 14478 16942 14530 16994
rect 17390 16942 17442 16994
rect 17614 16942 17666 16994
rect 20302 16942 20354 16994
rect 20638 16942 20690 16994
rect 24334 16942 24386 16994
rect 39230 16942 39282 16994
rect 40014 16942 40066 16994
rect 45054 16942 45106 16994
rect 49310 16942 49362 16994
rect 52894 16942 52946 16994
rect 1822 16830 1874 16882
rect 5070 16830 5122 16882
rect 6302 16830 6354 16882
rect 6526 16830 6578 16882
rect 7086 16830 7138 16882
rect 13134 16830 13186 16882
rect 13470 16830 13522 16882
rect 13582 16830 13634 16882
rect 14590 16830 14642 16882
rect 14814 16830 14866 16882
rect 15262 16830 15314 16882
rect 16046 16830 16098 16882
rect 16382 16830 16434 16882
rect 16606 16830 16658 16882
rect 17950 16830 18002 16882
rect 20078 16830 20130 16882
rect 20190 16830 20242 16882
rect 20974 16830 21026 16882
rect 23998 16830 24050 16882
rect 25230 16830 25282 16882
rect 36318 16830 36370 16882
rect 38558 16830 38610 16882
rect 38782 16830 38834 16882
rect 40238 16830 40290 16882
rect 43150 16830 43202 16882
rect 44494 16830 44546 16882
rect 49198 16830 49250 16882
rect 49534 16830 49586 16882
rect 52670 16830 52722 16882
rect 53230 16830 53282 16882
rect 4622 16718 4674 16770
rect 16158 16718 16210 16770
rect 17838 16718 17890 16770
rect 21646 16718 21698 16770
rect 23774 16718 23826 16770
rect 26014 16718 26066 16770
rect 28142 16718 28194 16770
rect 39230 16718 39282 16770
rect 42590 16718 42642 16770
rect 6862 16606 6914 16658
rect 14926 16606 14978 16658
rect 16494 16606 16546 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 15374 16270 15426 16322
rect 44718 16270 44770 16322
rect 44942 16270 44994 16322
rect 6078 16158 6130 16210
rect 12462 16158 12514 16210
rect 12798 16158 12850 16210
rect 17390 16158 17442 16210
rect 34862 16158 34914 16210
rect 42030 16158 42082 16210
rect 44270 16158 44322 16210
rect 44942 16158 44994 16210
rect 51214 16158 51266 16210
rect 4622 16046 4674 16098
rect 4958 16046 5010 16098
rect 6190 16046 6242 16098
rect 6862 16046 6914 16098
rect 9662 16046 9714 16098
rect 13582 16046 13634 16098
rect 15710 16046 15762 16098
rect 23102 16046 23154 16098
rect 23662 16046 23714 16098
rect 24446 16046 24498 16098
rect 25118 16046 25170 16098
rect 25678 16046 25730 16098
rect 34974 16046 35026 16098
rect 37550 16046 37602 16098
rect 39006 16046 39058 16098
rect 39454 16046 39506 16098
rect 40238 16046 40290 16098
rect 41246 16046 41298 16098
rect 42366 16046 42418 16098
rect 43822 16046 43874 16098
rect 48638 16046 48690 16098
rect 48862 16046 48914 16098
rect 49534 16046 49586 16098
rect 50094 16046 50146 16098
rect 50766 16046 50818 16098
rect 51886 16046 51938 16098
rect 52222 16046 52274 16098
rect 52894 16046 52946 16098
rect 53118 16046 53170 16098
rect 5070 15934 5122 15986
rect 6526 15934 6578 15986
rect 6638 15934 6690 15986
rect 10334 15934 10386 15986
rect 15486 15934 15538 15986
rect 17278 15934 17330 15986
rect 17502 15934 17554 15986
rect 23214 15934 23266 15986
rect 24670 15934 24722 15986
rect 25342 15934 25394 15986
rect 35646 15934 35698 15986
rect 38558 15934 38610 15986
rect 49198 15934 49250 15986
rect 49758 15934 49810 15986
rect 49982 15934 50034 15986
rect 50430 15934 50482 15986
rect 52670 15934 52722 15986
rect 12910 15822 12962 15874
rect 23326 15822 23378 15874
rect 23998 15822 24050 15874
rect 25566 15822 25618 15874
rect 37662 15822 37714 15874
rect 38446 15822 38498 15874
rect 48750 15822 48802 15874
rect 50654 15822 50706 15874
rect 51998 15822 52050 15874
rect 52782 15822 52834 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 6302 15486 6354 15538
rect 10446 15486 10498 15538
rect 18174 15486 18226 15538
rect 28814 15486 28866 15538
rect 34302 15486 34354 15538
rect 35310 15486 35362 15538
rect 39230 15486 39282 15538
rect 40238 15486 40290 15538
rect 41022 15486 41074 15538
rect 45502 15486 45554 15538
rect 46510 15486 46562 15538
rect 52334 15486 52386 15538
rect 5966 15374 6018 15426
rect 6078 15374 6130 15426
rect 8654 15374 8706 15426
rect 10334 15374 10386 15426
rect 10558 15374 10610 15426
rect 13582 15374 13634 15426
rect 13918 15374 13970 15426
rect 14254 15374 14306 15426
rect 14590 15374 14642 15426
rect 17390 15374 17442 15426
rect 17614 15374 17666 15426
rect 19518 15374 19570 15426
rect 33406 15374 33458 15426
rect 33966 15374 34018 15426
rect 36430 15374 36482 15426
rect 38782 15374 38834 15426
rect 48750 15374 48802 15426
rect 51774 15374 51826 15426
rect 8430 15262 8482 15314
rect 11118 15262 11170 15314
rect 17950 15262 18002 15314
rect 18846 15262 18898 15314
rect 22094 15262 22146 15314
rect 28478 15262 28530 15314
rect 29150 15262 29202 15314
rect 29598 15262 29650 15314
rect 36094 15262 36146 15314
rect 37326 15262 37378 15314
rect 39342 15262 39394 15314
rect 44158 15262 44210 15314
rect 44718 15262 44770 15314
rect 45838 15262 45890 15314
rect 46286 15262 46338 15314
rect 49086 15262 49138 15314
rect 51102 15262 51154 15314
rect 51438 15262 51490 15314
rect 21646 15150 21698 15202
rect 30382 15150 30434 15202
rect 32510 15150 32562 15202
rect 33518 15150 33570 15202
rect 41358 15150 41410 15202
rect 43486 15150 43538 15202
rect 48862 15150 48914 15202
rect 51326 15150 51378 15202
rect 52110 15150 52162 15202
rect 52222 15150 52274 15202
rect 10894 15038 10946 15090
rect 17838 15038 17890 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 6414 14702 6466 14754
rect 6638 14702 6690 14754
rect 36094 14702 36146 14754
rect 42254 14702 42306 14754
rect 9662 14590 9714 14642
rect 29374 14590 29426 14642
rect 31166 14590 31218 14642
rect 40798 14590 40850 14642
rect 42702 14590 42754 14642
rect 45838 14590 45890 14642
rect 48862 14590 48914 14642
rect 50990 14590 51042 14642
rect 52670 14590 52722 14642
rect 6190 14478 6242 14530
rect 8094 14478 8146 14530
rect 8318 14478 8370 14530
rect 8654 14478 8706 14530
rect 8878 14478 8930 14530
rect 9214 14478 9266 14530
rect 15150 14478 15202 14530
rect 15710 14478 15762 14530
rect 17390 14478 17442 14530
rect 17614 14478 17666 14530
rect 17726 14478 17778 14530
rect 19070 14478 19122 14530
rect 24334 14478 24386 14530
rect 26014 14478 26066 14530
rect 31502 14478 31554 14530
rect 31838 14478 31890 14530
rect 32062 14478 32114 14530
rect 39230 14478 39282 14530
rect 39790 14478 39842 14530
rect 42254 14478 42306 14530
rect 45390 14478 45442 14530
rect 46286 14478 46338 14530
rect 48190 14478 48242 14530
rect 6750 14366 6802 14418
rect 15374 14366 15426 14418
rect 17166 14366 17218 14418
rect 18286 14366 18338 14418
rect 18398 14366 18450 14418
rect 32286 14366 32338 14418
rect 35982 14366 36034 14418
rect 38782 14366 38834 14418
rect 39678 14366 39730 14418
rect 41918 14366 41970 14418
rect 46958 14366 47010 14418
rect 8206 14254 8258 14306
rect 9102 14254 9154 14306
rect 16046 14254 16098 14306
rect 17950 14254 18002 14306
rect 18510 14254 18562 14306
rect 23998 14254 24050 14306
rect 24222 14254 24274 14306
rect 26126 14254 26178 14306
rect 26350 14254 26402 14306
rect 31502 14254 31554 14306
rect 46510 14254 46562 14306
rect 46846 14254 46898 14306
rect 47406 14254 47458 14306
rect 51438 14254 51490 14306
rect 53230 14254 53282 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 5854 13918 5906 13970
rect 7310 13918 7362 13970
rect 7422 13918 7474 13970
rect 9662 13918 9714 13970
rect 10110 13918 10162 13970
rect 12686 13918 12738 13970
rect 13134 13918 13186 13970
rect 40014 13918 40066 13970
rect 46398 13918 46450 13970
rect 53342 13918 53394 13970
rect 5294 13806 5346 13858
rect 7534 13806 7586 13858
rect 8766 13806 8818 13858
rect 8878 13806 8930 13858
rect 10446 13806 10498 13858
rect 10894 13806 10946 13858
rect 11230 13806 11282 13858
rect 11566 13806 11618 13858
rect 12350 13806 12402 13858
rect 20974 13806 21026 13858
rect 39342 13806 39394 13858
rect 40126 13806 40178 13858
rect 46734 13806 46786 13858
rect 1822 13694 1874 13746
rect 4958 13694 5010 13746
rect 5630 13694 5682 13746
rect 7982 13694 8034 13746
rect 8654 13694 8706 13746
rect 11902 13694 11954 13746
rect 24670 13694 24722 13746
rect 25790 13694 25842 13746
rect 26014 13694 26066 13746
rect 26350 13694 26402 13746
rect 26574 13694 26626 13746
rect 36094 13694 36146 13746
rect 36654 13694 36706 13746
rect 38558 13694 38610 13746
rect 39118 13694 39170 13746
rect 39678 13694 39730 13746
rect 39902 13694 39954 13746
rect 40238 13694 40290 13746
rect 44718 13694 44770 13746
rect 45166 13694 45218 13746
rect 2494 13582 2546 13634
rect 4622 13582 4674 13634
rect 11790 13582 11842 13634
rect 21758 13582 21810 13634
rect 23886 13582 23938 13634
rect 25342 13582 25394 13634
rect 26126 13582 26178 13634
rect 27358 13582 27410 13634
rect 29486 13582 29538 13634
rect 35758 13582 35810 13634
rect 41806 13582 41858 13634
rect 43934 13582 43986 13634
rect 5966 13470 6018 13522
rect 8206 13470 8258 13522
rect 20862 13470 20914 13522
rect 38670 13470 38722 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15934 13134 15986 13186
rect 17614 13134 17666 13186
rect 18286 13134 18338 13186
rect 37886 13134 37938 13186
rect 42590 13134 42642 13186
rect 10782 13022 10834 13074
rect 12238 13022 12290 13074
rect 14590 13022 14642 13074
rect 19070 13022 19122 13074
rect 24110 13022 24162 13074
rect 33630 13022 33682 13074
rect 35422 13022 35474 13074
rect 37550 13022 37602 13074
rect 41022 13022 41074 13074
rect 43038 13022 43090 13074
rect 2606 12910 2658 12962
rect 8542 12910 8594 12962
rect 11454 12910 11506 12962
rect 15598 12910 15650 12962
rect 16382 12910 16434 12962
rect 17166 12910 17218 12962
rect 17390 12910 17442 12962
rect 17838 12910 17890 12962
rect 18398 12910 18450 12962
rect 18622 12910 18674 12962
rect 26126 12910 26178 12962
rect 26350 12910 26402 12962
rect 26686 12910 26738 12962
rect 30718 12910 30770 12962
rect 35982 12910 36034 12962
rect 38222 12910 38274 12962
rect 38670 12910 38722 12962
rect 39118 12910 39170 12962
rect 40910 12910 40962 12962
rect 42254 12910 42306 12962
rect 2270 12798 2322 12850
rect 8430 12798 8482 12850
rect 13806 12798 13858 12850
rect 16158 12798 16210 12850
rect 16830 12798 16882 12850
rect 31502 12798 31554 12850
rect 34638 12798 34690 12850
rect 35534 12798 35586 12850
rect 35758 12798 35810 12850
rect 39566 12798 39618 12850
rect 40462 12798 40514 12850
rect 42478 12798 42530 12850
rect 4846 12686 4898 12738
rect 8206 12686 8258 12738
rect 11230 12686 11282 12738
rect 13470 12686 13522 12738
rect 15934 12686 15986 12738
rect 17614 12686 17666 12738
rect 26574 12686 26626 12738
rect 27134 12686 27186 12738
rect 34302 12686 34354 12738
rect 36430 12686 36482 12738
rect 37998 12686 38050 12738
rect 40686 12686 40738 12738
rect 41022 12686 41074 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 7758 12350 7810 12402
rect 7870 12350 7922 12402
rect 8430 12350 8482 12402
rect 15150 12350 15202 12402
rect 19966 12350 20018 12402
rect 23886 12350 23938 12402
rect 28254 12350 28306 12402
rect 31838 12350 31890 12402
rect 35086 12350 35138 12402
rect 35310 12350 35362 12402
rect 35422 12350 35474 12402
rect 36094 12350 36146 12402
rect 36206 12350 36258 12402
rect 38670 12350 38722 12402
rect 44606 12350 44658 12402
rect 44942 12350 44994 12402
rect 46062 12350 46114 12402
rect 49870 12350 49922 12402
rect 5966 12238 6018 12290
rect 7086 12238 7138 12290
rect 14142 12238 14194 12290
rect 14366 12238 14418 12290
rect 14926 12238 14978 12290
rect 17390 12238 17442 12290
rect 23550 12238 23602 12290
rect 24110 12238 24162 12290
rect 24558 12238 24610 12290
rect 36318 12238 36370 12290
rect 39006 12238 39058 12290
rect 51102 12238 51154 12290
rect 5518 12126 5570 12178
rect 6414 12126 6466 12178
rect 6638 12126 6690 12178
rect 6862 12126 6914 12178
rect 7422 12126 7474 12178
rect 13582 12126 13634 12178
rect 13918 12126 13970 12178
rect 15598 12126 15650 12178
rect 15822 12126 15874 12178
rect 16046 12126 16098 12178
rect 16382 12126 16434 12178
rect 17614 12126 17666 12178
rect 17838 12126 17890 12178
rect 18062 12126 18114 12178
rect 23774 12126 23826 12178
rect 24334 12126 24386 12178
rect 24670 12126 24722 12178
rect 25790 12126 25842 12178
rect 32062 12126 32114 12178
rect 34750 12126 34802 12178
rect 35870 12126 35922 12178
rect 35982 12126 36034 12178
rect 38110 12126 38162 12178
rect 38334 12126 38386 12178
rect 44830 12126 44882 12178
rect 45054 12126 45106 12178
rect 49534 12126 49586 12178
rect 50318 12126 50370 12178
rect 5406 12014 5458 12066
rect 6078 12014 6130 12066
rect 6526 12014 6578 12066
rect 14254 12014 14306 12066
rect 15262 12014 15314 12066
rect 15710 12014 15762 12066
rect 17502 12014 17554 12066
rect 20414 12014 20466 12066
rect 26910 12014 26962 12066
rect 49198 12014 49250 12066
rect 53230 12014 53282 12066
rect 5182 11902 5234 11954
rect 7646 11902 7698 11954
rect 31726 11902 31778 11954
rect 37774 11902 37826 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6190 11566 6242 11618
rect 9102 11566 9154 11618
rect 9326 11566 9378 11618
rect 11118 11566 11170 11618
rect 13694 11566 13746 11618
rect 23214 11566 23266 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 6414 11454 6466 11506
rect 15822 11454 15874 11506
rect 17726 11454 17778 11506
rect 21422 11454 21474 11506
rect 27918 11454 27970 11506
rect 31726 11454 31778 11506
rect 32510 11454 32562 11506
rect 49086 11454 49138 11506
rect 1822 11342 1874 11394
rect 5742 11342 5794 11394
rect 8878 11342 8930 11394
rect 11454 11342 11506 11394
rect 12798 11342 12850 11394
rect 13470 11342 13522 11394
rect 14030 11342 14082 11394
rect 15262 11342 15314 11394
rect 20414 11342 20466 11394
rect 26574 11342 26626 11394
rect 27022 11342 27074 11394
rect 27358 11342 27410 11394
rect 29262 11342 29314 11394
rect 29486 11342 29538 11394
rect 30942 11342 30994 11394
rect 31166 11342 31218 11394
rect 31614 11342 31666 11394
rect 32174 11342 32226 11394
rect 32622 11342 32674 11394
rect 32846 11342 32898 11394
rect 40798 11342 40850 11394
rect 41470 11342 41522 11394
rect 45166 11342 45218 11394
rect 45838 11342 45890 11394
rect 46286 11342 46338 11394
rect 46958 11342 47010 11394
rect 5630 11230 5682 11282
rect 10670 11230 10722 11282
rect 10894 11230 10946 11282
rect 12910 11230 12962 11282
rect 14254 11230 14306 11282
rect 20750 11230 20802 11282
rect 23326 11230 23378 11282
rect 25902 11230 25954 11282
rect 26798 11230 26850 11282
rect 29150 11230 29202 11282
rect 45950 11230 46002 11282
rect 50654 11230 50706 11282
rect 52222 11230 52274 11282
rect 52894 11230 52946 11282
rect 53230 11230 53282 11282
rect 5070 11118 5122 11170
rect 6526 11118 6578 11170
rect 9774 11118 9826 11170
rect 11118 11118 11170 11170
rect 12686 11118 12738 11170
rect 13470 11118 13522 11170
rect 20638 11118 20690 11170
rect 23214 11118 23266 11170
rect 24334 11118 24386 11170
rect 26238 11118 26290 11170
rect 27358 11118 27410 11170
rect 31838 11118 31890 11170
rect 32398 11118 32450 11170
rect 41022 11118 41074 11170
rect 41694 11118 41746 11170
rect 42030 11118 42082 11170
rect 42366 11118 42418 11170
rect 42814 11118 42866 11170
rect 43262 11118 43314 11170
rect 45390 11118 45442 11170
rect 45614 11118 45666 11170
rect 49534 11118 49586 11170
rect 49982 11118 50034 11170
rect 50766 11118 50818 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 10334 10782 10386 10834
rect 17502 10782 17554 10834
rect 18734 10782 18786 10834
rect 19630 10782 19682 10834
rect 23774 10782 23826 10834
rect 23886 10782 23938 10834
rect 30382 10782 30434 10834
rect 30942 10782 30994 10834
rect 31950 10782 32002 10834
rect 32174 10782 32226 10834
rect 37326 10782 37378 10834
rect 40462 10782 40514 10834
rect 41358 10782 41410 10834
rect 41918 10782 41970 10834
rect 45614 10782 45666 10834
rect 49646 10782 49698 10834
rect 9550 10670 9602 10722
rect 9886 10670 9938 10722
rect 10558 10670 10610 10722
rect 11454 10670 11506 10722
rect 13694 10670 13746 10722
rect 13918 10670 13970 10722
rect 20750 10670 20802 10722
rect 23438 10670 23490 10722
rect 23550 10670 23602 10722
rect 24110 10670 24162 10722
rect 24222 10670 24274 10722
rect 25230 10670 25282 10722
rect 27582 10670 27634 10722
rect 31838 10670 31890 10722
rect 36430 10670 36482 10722
rect 36766 10670 36818 10722
rect 39006 10670 39058 10722
rect 39454 10670 39506 10722
rect 39566 10670 39618 10722
rect 42142 10670 42194 10722
rect 51102 10670 51154 10722
rect 5742 10558 5794 10610
rect 6078 10558 6130 10610
rect 6302 10558 6354 10610
rect 6638 10558 6690 10610
rect 7086 10558 7138 10610
rect 10110 10558 10162 10610
rect 10670 10558 10722 10610
rect 11118 10558 11170 10610
rect 16830 10558 16882 10610
rect 19966 10558 20018 10610
rect 25566 10558 25618 10610
rect 26910 10558 26962 10610
rect 30158 10558 30210 10610
rect 35646 10558 35698 10610
rect 35870 10558 35922 10610
rect 36206 10558 36258 10610
rect 38782 10558 38834 10610
rect 41134 10558 41186 10610
rect 41470 10558 41522 10610
rect 42926 10558 42978 10610
rect 43374 10558 43426 10610
rect 43822 10558 43874 10610
rect 45166 10558 45218 10610
rect 45390 10558 45442 10610
rect 49198 10558 49250 10610
rect 49422 10558 49474 10610
rect 49646 10558 49698 10610
rect 49870 10558 49922 10610
rect 50318 10558 50370 10610
rect 5630 10446 5682 10498
rect 6190 10446 6242 10498
rect 7422 10446 7474 10498
rect 9662 10446 9714 10498
rect 13582 10446 13634 10498
rect 15710 10446 15762 10498
rect 18846 10446 18898 10498
rect 22878 10446 22930 10498
rect 26014 10446 26066 10498
rect 29710 10446 29762 10498
rect 35982 10446 36034 10498
rect 41918 10446 41970 10498
rect 45054 10446 45106 10498
rect 53230 10446 53282 10498
rect 6526 10334 6578 10386
rect 39678 10334 39730 10386
rect 43934 10334 43986 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 11230 9998 11282 10050
rect 12462 9998 12514 10050
rect 14030 9998 14082 10050
rect 23550 9998 23602 10050
rect 27246 9998 27298 10050
rect 39230 9998 39282 10050
rect 44942 9998 44994 10050
rect 47406 9998 47458 10050
rect 2158 9886 2210 9938
rect 4286 9886 4338 9938
rect 10446 9886 10498 9938
rect 15038 9886 15090 9938
rect 17390 9886 17442 9938
rect 19518 9886 19570 9938
rect 29934 9886 29986 9938
rect 5070 9774 5122 9826
rect 11118 9774 11170 9826
rect 11566 9774 11618 9826
rect 11790 9774 11842 9826
rect 12350 9774 12402 9826
rect 12910 9774 12962 9826
rect 13918 9774 13970 9826
rect 14478 9774 14530 9826
rect 16606 9774 16658 9826
rect 23662 9774 23714 9826
rect 27134 9774 27186 9826
rect 29486 9774 29538 9826
rect 33854 9774 33906 9826
rect 36206 9774 36258 9826
rect 38446 9774 38498 9826
rect 38670 9774 38722 9826
rect 39118 9774 39170 9826
rect 41358 9774 41410 9826
rect 41806 9774 41858 9826
rect 45390 9774 45442 9826
rect 45614 9774 45666 9826
rect 45838 9774 45890 9826
rect 46398 9774 46450 9826
rect 46846 9774 46898 9826
rect 47854 9774 47906 9826
rect 48414 9774 48466 9826
rect 12686 9662 12738 9714
rect 14254 9662 14306 9714
rect 29150 9662 29202 9714
rect 36094 9662 36146 9714
rect 38894 9662 38946 9714
rect 40910 9662 40962 9714
rect 43598 9662 43650 9714
rect 46062 9662 46114 9714
rect 48078 9662 48130 9714
rect 48190 9662 48242 9714
rect 49534 9662 49586 9714
rect 49870 9662 49922 9714
rect 50206 9662 50258 9714
rect 50542 9662 50594 9714
rect 5742 9550 5794 9602
rect 11006 9550 11058 9602
rect 12126 9550 12178 9602
rect 14142 9550 14194 9602
rect 15374 9550 15426 9602
rect 16270 9550 16322 9602
rect 23550 9550 23602 9602
rect 27246 9550 27298 9602
rect 33630 9550 33682 9602
rect 35870 9550 35922 9602
rect 40798 9550 40850 9602
rect 46510 9550 46562 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 12126 9214 12178 9266
rect 13246 9214 13298 9266
rect 16718 9214 16770 9266
rect 26238 9214 26290 9266
rect 29822 9214 29874 9266
rect 31726 9214 31778 9266
rect 35646 9214 35698 9266
rect 36430 9214 36482 9266
rect 38334 9214 38386 9266
rect 42254 9214 42306 9266
rect 43822 9214 43874 9266
rect 23438 9102 23490 9154
rect 23774 9102 23826 9154
rect 31950 9102 32002 9154
rect 32174 9102 32226 9154
rect 33406 9102 33458 9154
rect 35870 9102 35922 9154
rect 36878 9102 36930 9154
rect 38110 9102 38162 9154
rect 29262 8990 29314 9042
rect 31054 8990 31106 9042
rect 31390 8990 31442 9042
rect 33070 8990 33122 9042
rect 35198 8990 35250 9042
rect 35422 8990 35474 9042
rect 36318 8990 36370 9042
rect 36654 8990 36706 9042
rect 42142 8990 42194 9042
rect 42478 8990 42530 9042
rect 45166 8990 45218 9042
rect 45390 8990 45442 9042
rect 45838 8990 45890 9042
rect 52222 8990 52274 9042
rect 52782 8990 52834 9042
rect 16830 8878 16882 8930
rect 26126 8878 26178 8930
rect 35310 8878 35362 8930
rect 38446 8878 38498 8930
rect 42814 8878 42866 8930
rect 45726 8878 45778 8930
rect 31726 8766 31778 8818
rect 33070 8766 33122 8818
rect 36766 8766 36818 8818
rect 45950 8766 46002 8818
rect 52558 8766 52610 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 12798 8430 12850 8482
rect 47294 8430 47346 8482
rect 8094 8318 8146 8370
rect 10222 8318 10274 8370
rect 15374 8318 15426 8370
rect 17502 8318 17554 8370
rect 22990 8318 23042 8370
rect 25342 8318 25394 8370
rect 26238 8318 26290 8370
rect 27246 8318 27298 8370
rect 31614 8318 31666 8370
rect 33742 8318 33794 8370
rect 36318 8318 36370 8370
rect 39342 8318 39394 8370
rect 7422 8206 7474 8258
rect 14590 8206 14642 8258
rect 19742 8206 19794 8258
rect 20302 8206 20354 8258
rect 20638 8206 20690 8258
rect 25230 8206 25282 8258
rect 25454 8206 25506 8258
rect 26014 8206 26066 8258
rect 26686 8206 26738 8258
rect 30830 8206 30882 8258
rect 35646 8206 35698 8258
rect 35870 8206 35922 8258
rect 37214 8206 37266 8258
rect 38894 8206 38946 8258
rect 41470 8206 41522 8258
rect 42702 8206 42754 8258
rect 42926 8206 42978 8258
rect 43150 8206 43202 8258
rect 43934 8206 43986 8258
rect 47182 8206 47234 8258
rect 49086 8206 49138 8258
rect 53230 8206 53282 8258
rect 12910 8094 12962 8146
rect 23550 8094 23602 8146
rect 24782 8094 24834 8146
rect 25790 8094 25842 8146
rect 26462 8094 26514 8146
rect 34750 8094 34802 8146
rect 34974 8094 35026 8146
rect 35422 8094 35474 8146
rect 35758 8094 35810 8146
rect 36990 8094 37042 8146
rect 39454 8094 39506 8146
rect 41806 8094 41858 8146
rect 43374 8094 43426 8146
rect 48638 8094 48690 8146
rect 49758 8094 49810 8146
rect 52894 8094 52946 8146
rect 10670 7982 10722 8034
rect 17950 7982 18002 8034
rect 19518 7982 19570 8034
rect 20526 7982 20578 8034
rect 22990 7982 23042 8034
rect 23102 7982 23154 8034
rect 23326 7982 23378 8034
rect 25006 7982 25058 8034
rect 26350 7982 26402 8034
rect 34862 7982 34914 8034
rect 39230 7982 39282 8034
rect 42590 7982 42642 8034
rect 43710 7982 43762 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 23102 7646 23154 7698
rect 23326 7646 23378 7698
rect 25902 7646 25954 7698
rect 31166 7646 31218 7698
rect 31838 7646 31890 7698
rect 39006 7646 39058 7698
rect 40910 7646 40962 7698
rect 42142 7646 42194 7698
rect 43710 7646 43762 7698
rect 46734 7646 46786 7698
rect 47070 7646 47122 7698
rect 53342 7646 53394 7698
rect 6078 7534 6130 7586
rect 11006 7534 11058 7586
rect 18510 7534 18562 7586
rect 20414 7534 20466 7586
rect 23550 7534 23602 7586
rect 28702 7534 28754 7586
rect 36094 7534 36146 7586
rect 36318 7534 36370 7586
rect 37886 7534 37938 7586
rect 38222 7534 38274 7586
rect 38334 7534 38386 7586
rect 38670 7534 38722 7586
rect 39566 7534 39618 7586
rect 42478 7534 42530 7586
rect 52334 7534 52386 7586
rect 5406 7422 5458 7474
rect 10222 7422 10274 7474
rect 18734 7422 18786 7474
rect 19630 7422 19682 7474
rect 22990 7422 23042 7474
rect 23214 7422 23266 7474
rect 26238 7422 26290 7474
rect 29486 7422 29538 7474
rect 36654 7422 36706 7474
rect 36990 7422 37042 7474
rect 37998 7422 38050 7474
rect 38894 7422 38946 7474
rect 39342 7422 39394 7474
rect 39790 7422 39842 7474
rect 41246 7422 41298 7474
rect 41694 7422 41746 7474
rect 46846 7422 46898 7474
rect 47742 7422 47794 7474
rect 47966 7422 48018 7474
rect 50094 7422 50146 7474
rect 52670 7422 52722 7474
rect 3502 7310 3554 7362
rect 8206 7310 8258 7362
rect 8542 7310 8594 7362
rect 13134 7310 13186 7362
rect 13582 7310 13634 7362
rect 16606 7310 16658 7362
rect 19294 7310 19346 7362
rect 22542 7310 22594 7362
rect 25454 7310 25506 7362
rect 26574 7310 26626 7362
rect 31054 7310 31106 7362
rect 36766 7310 36818 7362
rect 43038 7310 43090 7362
rect 49422 7310 49474 7362
rect 50206 7310 50258 7362
rect 3614 7198 3666 7250
rect 8654 7198 8706 7250
rect 8878 7198 8930 7250
rect 9102 7198 9154 7250
rect 18398 7198 18450 7250
rect 30942 7198 30994 7250
rect 41022 7198 41074 7250
rect 41806 7198 41858 7250
rect 46734 7198 46786 7250
rect 47518 7198 47570 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 32846 6862 32898 6914
rect 39230 6862 39282 6914
rect 43822 6862 43874 6914
rect 49982 6862 50034 6914
rect 16382 6750 16434 6802
rect 19854 6750 19906 6802
rect 45390 6750 45442 6802
rect 48526 6750 48578 6802
rect 8430 6638 8482 6690
rect 8878 6638 8930 6690
rect 9438 6638 9490 6690
rect 9662 6638 9714 6690
rect 13470 6638 13522 6690
rect 14254 6638 14306 6690
rect 17054 6638 17106 6690
rect 17726 6638 17778 6690
rect 27022 6638 27074 6690
rect 30718 6638 30770 6690
rect 33518 6638 33570 6690
rect 39118 6638 39170 6690
rect 40798 6638 40850 6690
rect 43374 6638 43426 6690
rect 43598 6638 43650 6690
rect 44046 6638 44098 6690
rect 44830 6638 44882 6690
rect 45726 6638 45778 6690
rect 46510 6638 46562 6690
rect 47406 6638 47458 6690
rect 47630 6638 47682 6690
rect 47854 6638 47906 6690
rect 48078 6638 48130 6690
rect 48414 6638 48466 6690
rect 49758 6638 49810 6690
rect 50206 6638 50258 6690
rect 50430 6638 50482 6690
rect 52670 6638 52722 6690
rect 9998 6526 10050 6578
rect 23886 6526 23938 6578
rect 31390 6526 31442 6578
rect 33406 6526 33458 6578
rect 40910 6526 40962 6578
rect 44270 6526 44322 6578
rect 46286 6526 46338 6578
rect 47182 6526 47234 6578
rect 48862 6526 48914 6578
rect 49534 6526 49586 6578
rect 50766 6526 50818 6578
rect 8990 6414 9042 6466
rect 9102 6414 9154 6466
rect 9886 6414 9938 6466
rect 10558 6414 10610 6466
rect 24222 6414 24274 6466
rect 26686 6414 26738 6466
rect 30382 6414 30434 6466
rect 31054 6414 31106 6466
rect 32510 6414 32562 6466
rect 34190 6414 34242 6466
rect 39230 6414 39282 6466
rect 41134 6414 41186 6466
rect 44382 6414 44434 6466
rect 47630 6414 47682 6466
rect 48638 6414 48690 6466
rect 50542 6414 50594 6466
rect 50878 6414 50930 6466
rect 52222 6414 52274 6466
rect 53230 6414 53282 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 9662 6078 9714 6130
rect 10334 6078 10386 6130
rect 14702 6078 14754 6130
rect 16606 6078 16658 6130
rect 22318 6078 22370 6130
rect 24110 6078 24162 6130
rect 24222 6078 24274 6130
rect 24446 6078 24498 6130
rect 27470 6078 27522 6130
rect 27806 6078 27858 6130
rect 9550 5966 9602 6018
rect 14814 5966 14866 6018
rect 22542 5966 22594 6018
rect 22766 5966 22818 6018
rect 34750 5966 34802 6018
rect 51102 5966 51154 6018
rect 22206 5854 22258 5906
rect 24558 5854 24610 5906
rect 27358 5854 27410 5906
rect 27694 5854 27746 5906
rect 33966 5854 34018 5906
rect 48750 5854 48802 5906
rect 49198 5854 49250 5906
rect 50318 5854 50370 5906
rect 22430 5742 22482 5794
rect 24334 5742 24386 5794
rect 27582 5742 27634 5794
rect 36878 5742 36930 5794
rect 37326 5742 37378 5794
rect 49982 5742 50034 5794
rect 53230 5742 53282 5794
rect 9662 5630 9714 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19518 5294 19570 5346
rect 25006 5294 25058 5346
rect 25342 5294 25394 5346
rect 28142 5294 28194 5346
rect 9774 5182 9826 5234
rect 11902 5182 11954 5234
rect 12350 5182 12402 5234
rect 15598 5182 15650 5234
rect 18846 5182 18898 5234
rect 19182 5182 19234 5234
rect 21310 5182 21362 5234
rect 22430 5182 22482 5234
rect 34078 5182 34130 5234
rect 38782 5182 38834 5234
rect 40910 5182 40962 5234
rect 44942 5182 44994 5234
rect 49534 5182 49586 5234
rect 8990 5070 9042 5122
rect 16046 5070 16098 5122
rect 16718 5070 16770 5122
rect 21646 5070 21698 5122
rect 22318 5070 22370 5122
rect 22542 5070 22594 5122
rect 22766 5070 22818 5122
rect 22990 5070 23042 5122
rect 25342 5070 25394 5122
rect 25790 5070 25842 5122
rect 27806 5070 27858 5122
rect 28478 5070 28530 5122
rect 31166 5070 31218 5122
rect 37998 5070 38050 5122
rect 46734 5070 46786 5122
rect 49982 5070 50034 5122
rect 31950 4958 32002 5010
rect 47406 4958 47458 5010
rect 19294 4846 19346 4898
rect 21422 4846 21474 4898
rect 28254 4846 28306 4898
rect 41358 4846 41410 4898
rect 44830 4846 44882 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 14926 4510 14978 4562
rect 31950 4510 32002 4562
rect 44494 4510 44546 4562
rect 47518 4510 47570 4562
rect 48862 4510 48914 4562
rect 49422 4510 49474 4562
rect 20750 4398 20802 4450
rect 25342 4398 25394 4450
rect 29934 4398 29986 4450
rect 32286 4398 32338 4450
rect 36206 4398 36258 4450
rect 41918 4398 41970 4450
rect 47630 4398 47682 4450
rect 49646 4398 49698 4450
rect 49982 4398 50034 4450
rect 51102 4398 51154 4450
rect 14366 4286 14418 4338
rect 19630 4286 19682 4338
rect 19966 4286 20018 4338
rect 30606 4286 30658 4338
rect 35422 4286 35474 4338
rect 38782 4286 38834 4338
rect 41246 4286 41298 4338
rect 50318 4286 50370 4338
rect 22878 4174 22930 4226
rect 27806 4174 27858 4226
rect 38334 4174 38386 4226
rect 44046 4174 44098 4226
rect 48078 4174 48130 4226
rect 53230 4174 53282 4226
rect 12126 4062 12178 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25342 3614 25394 3666
rect 27470 3614 27522 3666
rect 29822 3614 29874 3666
rect 36990 3614 37042 3666
rect 40238 3614 40290 3666
rect 42030 3614 42082 3666
rect 44382 3614 44434 3666
rect 46510 3614 46562 3666
rect 49646 3614 49698 3666
rect 52670 3614 52722 3666
rect 11902 3502 11954 3554
rect 24670 3502 24722 3554
rect 35534 3502 35586 3554
rect 35982 3502 36034 3554
rect 43710 3502 43762 3554
rect 47742 3502 47794 3554
rect 50654 3502 50706 3554
rect 2718 3390 2770 3442
rect 2942 3390 2994 3442
rect 3278 3390 3330 3442
rect 10110 3390 10162 3442
rect 12462 3390 12514 3442
rect 39342 3390 39394 3442
rect 39790 3390 39842 3442
rect 42478 3390 42530 3442
rect 42702 3390 42754 3442
rect 43038 3390 43090 3442
rect 47406 3390 47458 3442
rect 52446 3390 52498 3442
rect 53230 3390 53282 3442
rect 16942 3278 16994 3330
rect 20862 3278 20914 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 13664 54200 13776 55000
rect 41216 54200 41328 55000
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 13692 49028 13748 54200
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 41244 51604 41300 54200
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 41468 51604 41524 51614
rect 41244 51602 41524 51604
rect 41244 51550 41246 51602
rect 41298 51550 41470 51602
rect 41522 51550 41524 51602
rect 41244 51548 41524 51550
rect 41244 51538 41300 51548
rect 41468 51538 41524 51548
rect 51100 51604 51156 51614
rect 49868 51380 49924 51390
rect 32396 51266 32452 51278
rect 41916 51268 41972 51278
rect 32396 51214 32398 51266
rect 32450 51214 32452 51266
rect 19740 50708 19796 50718
rect 19628 50706 19796 50708
rect 19628 50654 19742 50706
rect 19794 50654 19796 50706
rect 19628 50652 19796 50654
rect 16940 50596 16996 50606
rect 16940 50502 16996 50540
rect 17948 50596 18004 50606
rect 17612 50484 17668 50494
rect 17612 50390 17668 50428
rect 13692 48972 13860 49028
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 12572 47570 12628 47582
rect 12572 47518 12574 47570
rect 12626 47518 12628 47570
rect 9772 47458 9828 47470
rect 9772 47406 9774 47458
rect 9826 47406 9828 47458
rect 9324 47236 9380 47246
rect 9772 47236 9828 47406
rect 10444 47348 10500 47358
rect 10444 47346 10948 47348
rect 10444 47294 10446 47346
rect 10498 47294 10948 47346
rect 10444 47292 10948 47294
rect 10444 47282 10500 47292
rect 9324 47234 9828 47236
rect 9324 47182 9326 47234
rect 9378 47182 9828 47234
rect 9324 47180 9828 47182
rect 9324 47170 9380 47180
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 7308 45444 7364 45454
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 6860 44324 6916 44334
rect 7308 44324 7364 45388
rect 9772 45444 9828 47180
rect 10892 46002 10948 47292
rect 10892 45950 10894 46002
rect 10946 45950 10948 46002
rect 10892 45938 10948 45950
rect 10780 45890 10836 45902
rect 10780 45838 10782 45890
rect 10834 45838 10836 45890
rect 10444 45780 10500 45790
rect 10332 45724 10444 45780
rect 9828 45388 10164 45444
rect 9772 45350 9828 45388
rect 9660 44436 9716 44446
rect 9660 44342 9716 44380
rect 10108 44434 10164 45388
rect 10108 44382 10110 44434
rect 10162 44382 10164 44434
rect 10108 44370 10164 44382
rect 6860 44322 7364 44324
rect 6860 44270 6862 44322
rect 6914 44270 7364 44322
rect 6860 44268 7364 44270
rect 6860 44258 6916 44268
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 7308 41186 7364 44268
rect 7532 44210 7588 44222
rect 7532 44158 7534 44210
rect 7586 44158 7588 44210
rect 7532 43652 7588 44158
rect 7532 43586 7588 43596
rect 9660 44100 9716 44110
rect 9660 43650 9716 44044
rect 9996 43876 10052 43886
rect 9660 43598 9662 43650
rect 9714 43598 9716 43650
rect 9660 43586 9716 43598
rect 9772 43652 9828 43662
rect 9772 43558 9828 43596
rect 9996 43650 10052 43820
rect 9996 43598 9998 43650
rect 10050 43598 10052 43650
rect 9996 43586 10052 43598
rect 10220 43540 10276 43550
rect 10332 43540 10388 45724
rect 10444 45686 10500 45724
rect 10780 45444 10836 45838
rect 11116 45890 11172 45902
rect 11116 45838 11118 45890
rect 11170 45838 11172 45890
rect 10780 45388 11060 45444
rect 11004 45330 11060 45388
rect 11004 45278 11006 45330
rect 11058 45278 11060 45330
rect 11004 45266 11060 45278
rect 11116 45332 11172 45838
rect 11228 45780 11284 45790
rect 11452 45780 11508 45790
rect 11284 45778 11508 45780
rect 11284 45726 11454 45778
rect 11506 45726 11508 45778
rect 11284 45724 11508 45726
rect 11228 45714 11284 45724
rect 11452 45714 11508 45724
rect 11116 45266 11172 45276
rect 12348 45332 12404 45342
rect 12236 45220 12292 45230
rect 12236 45126 12292 45164
rect 10892 45106 10948 45118
rect 11116 45108 11172 45118
rect 10892 45054 10894 45106
rect 10946 45054 10948 45106
rect 10892 44548 10948 45054
rect 10668 44492 10892 44548
rect 10444 44436 10500 44446
rect 10500 44380 10612 44436
rect 10444 44370 10500 44380
rect 10556 43708 10612 44380
rect 10668 44322 10724 44492
rect 10892 44482 10948 44492
rect 11004 45106 11172 45108
rect 11004 45054 11118 45106
rect 11170 45054 11172 45106
rect 11004 45052 11172 45054
rect 10668 44270 10670 44322
rect 10722 44270 10724 44322
rect 10668 44258 10724 44270
rect 10780 44100 10836 44110
rect 10780 44006 10836 44044
rect 10892 44100 10948 44110
rect 11004 44100 11060 45052
rect 11116 45042 11172 45052
rect 11564 45106 11620 45118
rect 11564 45054 11566 45106
rect 11618 45054 11620 45106
rect 11564 44996 11620 45054
rect 11564 44930 11620 44940
rect 11788 45106 11844 45118
rect 11788 45054 11790 45106
rect 11842 45054 11844 45106
rect 11788 44772 11844 45054
rect 12012 45106 12068 45118
rect 12012 45054 12014 45106
rect 12066 45054 12068 45106
rect 11676 44716 11956 44772
rect 11340 44324 11396 44334
rect 10892 44098 11060 44100
rect 10892 44046 10894 44098
rect 10946 44046 11060 44098
rect 10892 44044 11060 44046
rect 11116 44268 11340 44324
rect 10892 43988 10948 44044
rect 10892 43922 10948 43932
rect 11116 43762 11172 44268
rect 11340 44230 11396 44268
rect 11676 44210 11732 44716
rect 11788 44548 11844 44558
rect 11788 44322 11844 44492
rect 11900 44436 11956 44716
rect 11900 44370 11956 44380
rect 11788 44270 11790 44322
rect 11842 44270 11844 44322
rect 11788 44258 11844 44270
rect 11676 44158 11678 44210
rect 11730 44158 11732 44210
rect 11676 44146 11732 44158
rect 11452 44098 11508 44110
rect 11452 44046 11454 44098
rect 11506 44046 11508 44098
rect 11452 43876 11508 44046
rect 11452 43810 11508 43820
rect 12012 43876 12068 45054
rect 12348 44882 12404 45276
rect 12460 45108 12516 45118
rect 12460 45014 12516 45052
rect 12572 44996 12628 47518
rect 13020 47460 13076 47470
rect 13020 46674 13076 47404
rect 13020 46622 13022 46674
rect 13074 46622 13076 46674
rect 13020 46610 13076 46622
rect 13692 46564 13748 46574
rect 13692 46470 13748 46508
rect 12572 44930 12628 44940
rect 12684 45220 12740 45230
rect 12348 44830 12350 44882
rect 12402 44830 12404 44882
rect 12348 44818 12404 44830
rect 12572 44436 12628 44446
rect 12572 44322 12628 44380
rect 12572 44270 12574 44322
rect 12626 44270 12628 44322
rect 12572 44258 12628 44270
rect 12684 44324 12740 45164
rect 12908 45220 12964 45230
rect 12908 45126 12964 45164
rect 13356 45106 13412 45118
rect 13356 45054 13358 45106
rect 13410 45054 13412 45106
rect 12908 44994 12964 45006
rect 12908 44942 12910 44994
rect 12962 44942 12964 44994
rect 12684 44230 12740 44268
rect 12796 44884 12852 44894
rect 12796 44322 12852 44828
rect 12908 44548 12964 44942
rect 12908 44482 12964 44492
rect 13356 44436 13412 45054
rect 13356 44370 13412 44380
rect 12796 44270 12798 44322
rect 12850 44270 12852 44322
rect 12796 44212 12852 44270
rect 12796 44146 12852 44156
rect 13580 44212 13636 44222
rect 11116 43710 11118 43762
rect 11170 43710 11172 43762
rect 10556 43652 10948 43708
rect 11116 43698 11172 43710
rect 10220 43538 10388 43540
rect 10220 43486 10222 43538
rect 10274 43486 10388 43538
rect 10220 43484 10388 43486
rect 10220 43474 10276 43484
rect 10332 42532 10388 43484
rect 10892 43540 10948 43652
rect 10892 43446 10948 43484
rect 11788 43540 11844 43550
rect 10444 42532 10500 42542
rect 10892 42532 10948 42542
rect 10332 42530 10948 42532
rect 10332 42478 10446 42530
rect 10498 42478 10894 42530
rect 10946 42478 10948 42530
rect 10332 42476 10948 42478
rect 10220 41972 10276 41982
rect 10332 41972 10388 42476
rect 10444 42466 10500 42476
rect 10892 42466 10948 42476
rect 11676 42196 11732 42206
rect 11228 42140 11676 42196
rect 10892 42082 10948 42094
rect 10892 42030 10894 42082
rect 10946 42030 10948 42082
rect 10220 41970 10388 41972
rect 10220 41918 10222 41970
rect 10274 41918 10388 41970
rect 10220 41916 10388 41918
rect 10220 41906 10276 41916
rect 8092 41860 8148 41870
rect 8092 41298 8148 41804
rect 8092 41246 8094 41298
rect 8146 41246 8148 41298
rect 8092 41234 8148 41246
rect 10220 41298 10276 41310
rect 10220 41246 10222 41298
rect 10274 41246 10276 41298
rect 7308 41134 7310 41186
rect 7362 41134 7364 41186
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5740 39620 5796 39630
rect 5740 39526 5796 39564
rect 7308 39620 7364 41134
rect 10220 41188 10276 41246
rect 10220 41122 10276 41132
rect 7308 39554 7364 39564
rect 8540 39730 8596 39742
rect 8540 39678 8542 39730
rect 8594 39678 8596 39730
rect 6412 39508 6468 39518
rect 6412 39506 6916 39508
rect 6412 39454 6414 39506
rect 6466 39454 6916 39506
rect 6412 39452 6916 39454
rect 6412 39442 6468 39452
rect 6860 39058 6916 39452
rect 6860 39006 6862 39058
rect 6914 39006 6916 39058
rect 6860 38994 6916 39006
rect 6524 38836 6580 38846
rect 6524 38668 6580 38780
rect 6412 38612 6580 38668
rect 6860 38834 6916 38846
rect 7084 38836 7140 38846
rect 6860 38782 6862 38834
rect 6914 38782 6916 38834
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5516 37436 5908 37492
rect 5180 37380 5236 37390
rect 5068 37378 5236 37380
rect 5068 37326 5182 37378
rect 5234 37326 5236 37378
rect 5068 37324 5236 37326
rect 1820 37266 1876 37278
rect 1820 37214 1822 37266
rect 1874 37214 1876 37266
rect 1820 35028 1876 37214
rect 2492 37156 2548 37166
rect 2492 37062 2548 37100
rect 4620 37156 4676 37166
rect 5068 37156 5124 37324
rect 5180 37314 5236 37324
rect 5292 37268 5348 37278
rect 5292 37174 5348 37212
rect 4620 37154 5124 37156
rect 4620 37102 4622 37154
rect 4674 37102 5124 37154
rect 4620 37100 5124 37102
rect 4620 37090 4676 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36258 4900 36270
rect 4844 36206 4846 36258
rect 4898 36206 4900 36258
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1820 34914 1876 34972
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 34850 1876 34862
rect 4620 35026 4676 35038
rect 4620 34974 4622 35026
rect 4674 34974 4676 35026
rect 2492 34804 2548 34814
rect 2492 34710 2548 34748
rect 4620 34132 4676 34974
rect 4844 35028 4900 36206
rect 5068 35700 5124 37100
rect 5180 37044 5236 37054
rect 5516 37044 5572 37436
rect 5180 37042 5572 37044
rect 5180 36990 5182 37042
rect 5234 36990 5572 37042
rect 5180 36988 5572 36990
rect 5628 37266 5684 37278
rect 5628 37214 5630 37266
rect 5682 37214 5684 37266
rect 5180 36978 5236 36988
rect 5628 36708 5684 37214
rect 5852 37266 5908 37436
rect 5852 37214 5854 37266
rect 5906 37214 5908 37266
rect 5852 37202 5908 37214
rect 6188 37268 6244 37278
rect 6412 37268 6468 38612
rect 6860 38274 6916 38782
rect 6972 38834 7140 38836
rect 6972 38782 7086 38834
rect 7138 38782 7140 38834
rect 6972 38780 7140 38782
rect 6972 38668 7028 38780
rect 7084 38770 7140 38780
rect 6972 38612 7140 38668
rect 6860 38222 6862 38274
rect 6914 38222 6916 38274
rect 6860 38210 6916 38222
rect 6972 38052 7028 38062
rect 6748 38050 7028 38052
rect 6748 37998 6974 38050
rect 7026 37998 7028 38050
rect 6748 37996 7028 37998
rect 6188 37266 6468 37268
rect 6188 37214 6190 37266
rect 6242 37214 6468 37266
rect 6188 37212 6468 37214
rect 6188 37202 6244 37212
rect 5740 37156 5796 37166
rect 5740 37062 5796 37100
rect 5740 36708 5796 36718
rect 5628 36706 5796 36708
rect 5628 36654 5742 36706
rect 5794 36654 5796 36706
rect 5628 36652 5796 36654
rect 5740 36642 5796 36652
rect 5516 36484 5572 36494
rect 5292 36482 5572 36484
rect 5292 36430 5518 36482
rect 5570 36430 5572 36482
rect 5292 36428 5572 36430
rect 5292 35922 5348 36428
rect 5516 36418 5572 36428
rect 5852 36258 5908 36270
rect 5852 36206 5854 36258
rect 5906 36206 5908 36258
rect 5740 35924 5796 35934
rect 5292 35870 5294 35922
rect 5346 35870 5348 35922
rect 5292 35858 5348 35870
rect 5404 35868 5740 35924
rect 5068 35634 5124 35644
rect 5180 35810 5236 35822
rect 5180 35758 5182 35810
rect 5234 35758 5236 35810
rect 5180 35252 5236 35758
rect 5404 35810 5460 35868
rect 5740 35830 5796 35868
rect 5404 35758 5406 35810
rect 5458 35758 5460 35810
rect 5404 35746 5460 35758
rect 5852 35700 5908 36206
rect 6076 36260 6132 36270
rect 6300 36260 6356 36270
rect 6076 36258 6300 36260
rect 6076 36206 6078 36258
rect 6130 36206 6300 36258
rect 6076 36204 6300 36206
rect 6076 36194 6132 36204
rect 6300 35810 6356 36204
rect 6300 35758 6302 35810
rect 6354 35758 6356 35810
rect 6300 35746 6356 35758
rect 6188 35700 6244 35710
rect 5852 35698 6244 35700
rect 5852 35646 6190 35698
rect 6242 35646 6244 35698
rect 5852 35644 6244 35646
rect 5180 35196 5572 35252
rect 4844 34962 4900 34972
rect 5180 35028 5236 35038
rect 5180 34934 5236 34972
rect 4620 34066 4676 34076
rect 5292 34132 5348 34142
rect 5292 34038 5348 34076
rect 5516 33906 5572 35196
rect 6188 34468 6244 35644
rect 6412 35476 6468 37212
rect 6636 37266 6692 37278
rect 6636 37214 6638 37266
rect 6690 37214 6692 37266
rect 6636 36036 6692 37214
rect 6748 37268 6804 37996
rect 6972 37986 7028 37996
rect 6860 37828 6916 37838
rect 6860 37734 6916 37772
rect 7084 37716 7140 38612
rect 6972 37660 7140 37716
rect 7532 37828 7588 37838
rect 6748 36932 6804 37212
rect 6860 37266 6916 37278
rect 6860 37214 6862 37266
rect 6914 37214 6916 37266
rect 6860 37156 6916 37214
rect 6860 37090 6916 37100
rect 6972 37154 7028 37660
rect 7084 37380 7140 37390
rect 7420 37380 7476 37390
rect 7084 37378 7476 37380
rect 7084 37326 7086 37378
rect 7138 37326 7422 37378
rect 7474 37326 7476 37378
rect 7084 37324 7476 37326
rect 7084 37314 7140 37324
rect 7420 37314 7476 37324
rect 6972 37102 6974 37154
rect 7026 37102 7028 37154
rect 6972 37090 7028 37102
rect 7532 37156 7588 37772
rect 7532 37062 7588 37100
rect 8540 37156 8596 39678
rect 8540 37090 8596 37100
rect 8988 39732 9044 39742
rect 8988 37156 9044 39676
rect 10108 39618 10164 39630
rect 10108 39566 10110 39618
rect 10162 39566 10164 39618
rect 10108 39508 10164 39566
rect 10332 39620 10388 41916
rect 10444 41972 10500 41982
rect 10444 41878 10500 41916
rect 10780 41972 10836 41982
rect 10892 41972 10948 42030
rect 10780 41970 10948 41972
rect 10780 41918 10782 41970
rect 10834 41918 10948 41970
rect 10780 41916 10948 41918
rect 11116 42082 11172 42094
rect 11116 42030 11118 42082
rect 11170 42030 11172 42082
rect 10780 41906 10836 41916
rect 10556 41860 10612 41870
rect 10556 41766 10612 41804
rect 10892 41188 10948 41198
rect 10780 40628 10836 40638
rect 10780 40534 10836 40572
rect 10892 40404 10948 41132
rect 11116 41076 11172 42030
rect 11228 42082 11284 42140
rect 11676 42102 11732 42140
rect 11228 42030 11230 42082
rect 11282 42030 11284 42082
rect 11228 42018 11284 42030
rect 11116 40982 11172 41020
rect 11564 40962 11620 40974
rect 11564 40910 11566 40962
rect 11618 40910 11620 40962
rect 10892 40338 10948 40348
rect 11228 40628 11284 40638
rect 10556 39620 10612 39630
rect 10332 39618 10724 39620
rect 10332 39566 10558 39618
rect 10610 39566 10724 39618
rect 10332 39564 10724 39566
rect 10556 39554 10612 39564
rect 10108 39060 10164 39452
rect 10556 39060 10612 39070
rect 10108 39058 10612 39060
rect 10108 39006 10110 39058
rect 10162 39006 10558 39058
rect 10610 39006 10612 39058
rect 10108 39004 10612 39006
rect 10108 38994 10164 39004
rect 10556 38994 10612 39004
rect 9772 38948 9828 38958
rect 9772 38854 9828 38892
rect 10668 38836 10724 39564
rect 11004 39618 11060 39630
rect 11004 39566 11006 39618
rect 11058 39566 11060 39618
rect 11004 39060 11060 39566
rect 11228 39508 11284 40572
rect 11564 39732 11620 40910
rect 11564 39666 11620 39676
rect 11284 39452 11620 39508
rect 11228 39414 11284 39452
rect 11004 38994 11060 39004
rect 10668 38780 11172 38836
rect 9548 37266 9604 37278
rect 9548 37214 9550 37266
rect 9602 37214 9604 37266
rect 9548 37156 9604 37214
rect 8988 37154 9604 37156
rect 8988 37102 8990 37154
rect 9042 37102 9604 37154
rect 8988 37100 9604 37102
rect 9884 37156 9940 37166
rect 10332 37156 10388 37166
rect 6748 36876 7028 36932
rect 6636 35980 6916 36036
rect 6636 35924 6692 35980
rect 6636 35858 6692 35868
rect 6860 35922 6916 35980
rect 6860 35870 6862 35922
rect 6914 35870 6916 35922
rect 6860 35858 6916 35870
rect 6972 35922 7028 36876
rect 6972 35870 6974 35922
rect 7026 35870 7028 35922
rect 6972 35858 7028 35870
rect 7308 35810 7364 35822
rect 7308 35758 7310 35810
rect 7362 35758 7364 35810
rect 6524 35700 6580 35710
rect 6524 35606 6580 35644
rect 7084 35698 7140 35710
rect 7084 35646 7086 35698
rect 7138 35646 7140 35698
rect 6412 35420 6692 35476
rect 6188 34402 6244 34412
rect 6524 34804 6580 34814
rect 6524 34354 6580 34748
rect 6524 34302 6526 34354
rect 6578 34302 6580 34354
rect 6524 34290 6580 34302
rect 6188 34132 6244 34142
rect 6412 34132 6468 34142
rect 6188 34130 6468 34132
rect 6188 34078 6190 34130
rect 6242 34078 6414 34130
rect 6466 34078 6468 34130
rect 6188 34076 6468 34078
rect 6188 34066 6244 34076
rect 6412 34066 6468 34076
rect 6636 34020 6692 35420
rect 6748 34244 6804 34254
rect 6748 34150 6804 34188
rect 6972 34130 7028 34142
rect 6972 34078 6974 34130
rect 7026 34078 7028 34130
rect 6972 34020 7028 34078
rect 6636 33964 7028 34020
rect 5516 33854 5518 33906
rect 5570 33854 5572 33906
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1820 32562 1876 32574
rect 1820 32510 1822 32562
rect 1874 32510 1876 32562
rect 1820 32452 1876 32510
rect 4956 32564 5012 32574
rect 1820 31948 1876 32396
rect 1708 31892 1876 31948
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 31892 2548 32398
rect 4620 32450 4676 32462
rect 4620 32398 4622 32450
rect 4674 32398 4676 32450
rect 4620 32340 4676 32398
rect 4620 32284 4900 32340
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1708 30210 1764 31892
rect 2492 31826 2548 31836
rect 4732 31668 4788 31678
rect 4844 31668 4900 32284
rect 4956 31890 5012 32508
rect 4956 31838 4958 31890
rect 5010 31838 5012 31890
rect 4956 31826 5012 31838
rect 5180 32452 5236 32462
rect 5068 31778 5124 31790
rect 5068 31726 5070 31778
rect 5122 31726 5124 31778
rect 5068 31668 5124 31726
rect 4844 31612 5124 31668
rect 4732 31574 4788 31612
rect 5068 31556 5124 31612
rect 5068 31490 5124 31500
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4620 30324 4676 30334
rect 4620 30230 4676 30268
rect 1708 30158 1710 30210
rect 1762 30158 1764 30210
rect 1708 27858 1764 30158
rect 5068 30212 5124 30222
rect 5180 30212 5236 32396
rect 5068 30210 5236 30212
rect 5068 30158 5070 30210
rect 5122 30158 5236 30210
rect 5068 30156 5236 30158
rect 5292 31668 5348 31678
rect 5516 31668 5572 33854
rect 5740 33906 5796 33918
rect 5740 33854 5742 33906
rect 5794 33854 5796 33906
rect 5740 33460 5796 33854
rect 6972 33684 7028 33964
rect 6972 33618 7028 33628
rect 5740 33394 5796 33404
rect 5740 32674 5796 32686
rect 5740 32622 5742 32674
rect 5794 32622 5796 32674
rect 5628 32564 5684 32574
rect 5628 32470 5684 32508
rect 5740 31892 5796 32622
rect 5964 32562 6020 32574
rect 5964 32510 5966 32562
rect 6018 32510 6020 32562
rect 5348 31612 5572 31668
rect 5628 31836 5796 31892
rect 5852 31892 5908 31902
rect 2492 30100 2548 30110
rect 2492 30006 2548 30044
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4956 27860 5012 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 24722 1764 27806
rect 4620 27804 4956 27860
rect 2492 27748 2548 27758
rect 2492 27654 2548 27692
rect 4620 27746 4676 27804
rect 4956 27766 5012 27804
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27682 4676 27694
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 27188 4900 27198
rect 5068 27188 5124 30156
rect 5292 30100 5348 31612
rect 5628 30996 5684 31836
rect 5852 31798 5908 31836
rect 5964 31778 6020 32510
rect 6412 32452 6468 32462
rect 6412 32358 6468 32396
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31714 6020 31726
rect 6300 31892 6356 31902
rect 6300 31778 6356 31836
rect 6300 31726 6302 31778
rect 6354 31726 6356 31778
rect 6300 31714 6356 31726
rect 5740 31666 5796 31678
rect 5740 31614 5742 31666
rect 5794 31614 5796 31666
rect 5740 31332 5796 31614
rect 6860 31666 6916 31678
rect 6860 31614 6862 31666
rect 6914 31614 6916 31666
rect 6524 31556 6580 31566
rect 6412 31554 6580 31556
rect 6412 31502 6526 31554
rect 6578 31502 6580 31554
rect 6412 31500 6580 31502
rect 6412 31444 6468 31500
rect 6524 31490 6580 31500
rect 6748 31556 6804 31566
rect 6748 31462 6804 31500
rect 5964 31388 6468 31444
rect 5964 31332 6020 31388
rect 5740 31276 6020 31332
rect 6636 31220 6692 31230
rect 6860 31220 6916 31614
rect 6188 31218 6916 31220
rect 6188 31166 6638 31218
rect 6690 31166 6916 31218
rect 6188 31164 6916 31166
rect 6076 31106 6132 31118
rect 6076 31054 6078 31106
rect 6130 31054 6132 31106
rect 6076 30996 6132 31054
rect 6188 31106 6244 31164
rect 6636 31154 6692 31164
rect 6188 31054 6190 31106
rect 6242 31054 6244 31106
rect 6188 31042 6244 31054
rect 5628 30930 5684 30940
rect 5740 30940 6132 30996
rect 6300 30996 6356 31006
rect 6524 30996 6580 31006
rect 6748 30996 6804 31006
rect 6356 30994 6692 30996
rect 6356 30942 6526 30994
rect 6578 30942 6692 30994
rect 6356 30940 6692 30942
rect 4844 27186 5124 27188
rect 4844 27134 4846 27186
rect 4898 27134 5124 27186
rect 4844 27132 5124 27134
rect 4844 27122 4900 27132
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 22370 1764 24670
rect 2940 25284 2996 25294
rect 2492 24612 2548 24622
rect 2492 24610 2660 24612
rect 2492 24558 2494 24610
rect 2546 24558 2660 24610
rect 2492 24556 2660 24558
rect 2492 24546 2548 24556
rect 2604 24162 2660 24556
rect 2604 24110 2606 24162
rect 2658 24110 2660 24162
rect 2604 24098 2660 24110
rect 2940 24162 2996 25228
rect 5068 24946 5124 27132
rect 5180 30044 5348 30100
rect 5740 30324 5796 30940
rect 6300 30930 6356 30940
rect 6524 30930 6580 30940
rect 6076 30772 6132 30782
rect 6076 30770 6468 30772
rect 6076 30718 6078 30770
rect 6130 30718 6468 30770
rect 6076 30716 6468 30718
rect 6076 30706 6132 30716
rect 5180 26908 5236 30044
rect 5740 28644 5796 30268
rect 6412 30210 6468 30716
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 6188 30098 6244 30110
rect 6188 30046 6190 30098
rect 6242 30046 6244 30098
rect 5740 28550 5796 28588
rect 5852 29538 5908 29550
rect 5852 29486 5854 29538
rect 5906 29486 5908 29538
rect 5852 28530 5908 29486
rect 6076 29426 6132 29438
rect 6076 29374 6078 29426
rect 6130 29374 6132 29426
rect 5852 28478 5854 28530
rect 5906 28478 5908 28530
rect 5852 28420 5908 28478
rect 5292 28364 5908 28420
rect 5964 28530 6020 28542
rect 5964 28478 5966 28530
rect 6018 28478 6020 28530
rect 5292 28084 5348 28364
rect 5964 28308 6020 28478
rect 5292 27970 5348 28028
rect 5292 27918 5294 27970
rect 5346 27918 5348 27970
rect 5292 27188 5348 27918
rect 5628 28252 6020 28308
rect 5628 27412 5684 28252
rect 5964 28084 6020 28094
rect 5964 28026 6020 28028
rect 5964 27974 5966 28026
rect 6018 27974 6020 28026
rect 5964 27962 6020 27974
rect 6076 27972 6132 29374
rect 6188 29314 6244 30046
rect 6300 30100 6356 30110
rect 6300 30006 6356 30044
rect 6412 29428 6468 29438
rect 6412 29334 6468 29372
rect 6188 29262 6190 29314
rect 6242 29262 6244 29314
rect 6188 29250 6244 29262
rect 6636 29204 6692 30940
rect 6748 30994 7028 30996
rect 6748 30942 6750 30994
rect 6802 30942 7028 30994
rect 6748 30940 7028 30942
rect 6748 30930 6804 30940
rect 6972 30212 7028 30940
rect 6748 30100 6804 30110
rect 6748 30006 6804 30044
rect 6860 29652 6916 29662
rect 6860 29558 6916 29596
rect 6748 29428 6804 29438
rect 6748 29334 6804 29372
rect 6972 29204 7028 30156
rect 7084 29764 7140 35646
rect 7196 34244 7252 34254
rect 7196 34150 7252 34188
rect 7196 30996 7252 31006
rect 7308 30996 7364 35758
rect 8428 35028 8484 35038
rect 8428 34934 8484 34972
rect 8988 35028 9044 37100
rect 9548 36932 9604 36942
rect 9604 36876 9716 36932
rect 9548 36866 9604 36876
rect 9548 36370 9604 36382
rect 9548 36318 9550 36370
rect 9602 36318 9604 36370
rect 8988 34962 9044 34972
rect 9212 36260 9268 36270
rect 7532 34914 7588 34926
rect 7532 34862 7534 34914
rect 7586 34862 7588 34914
rect 7532 34692 7588 34862
rect 9212 34916 9268 36204
rect 9548 35812 9604 36318
rect 9548 35718 9604 35756
rect 9660 34916 9716 36876
rect 9884 35924 9940 37100
rect 9996 37154 10388 37156
rect 9996 37102 10334 37154
rect 10386 37102 10388 37154
rect 9996 37100 10388 37102
rect 9996 36594 10052 37100
rect 10332 37090 10388 37100
rect 9996 36542 9998 36594
rect 10050 36542 10052 36594
rect 9996 36530 10052 36542
rect 10220 36370 10276 36382
rect 10220 36318 10222 36370
rect 10274 36318 10276 36370
rect 9996 36260 10052 36270
rect 9996 36166 10052 36204
rect 9996 35924 10052 35934
rect 9884 35868 9996 35924
rect 9996 35830 10052 35868
rect 9772 35700 9828 35710
rect 9772 35606 9828 35644
rect 9996 35586 10052 35598
rect 9996 35534 9998 35586
rect 10050 35534 10052 35586
rect 9884 34916 9940 34926
rect 9212 34850 9268 34860
rect 9324 34914 9940 34916
rect 9324 34862 9886 34914
rect 9938 34862 9940 34914
rect 9324 34860 9940 34862
rect 7532 34626 7588 34636
rect 8092 34468 8148 34478
rect 7532 34356 7588 34366
rect 7420 34242 7476 34254
rect 7420 34190 7422 34242
rect 7474 34190 7476 34242
rect 7420 34132 7476 34190
rect 7532 34242 7588 34300
rect 7532 34190 7534 34242
rect 7586 34190 7588 34242
rect 7532 34178 7588 34190
rect 7868 34356 7924 34366
rect 7420 34066 7476 34076
rect 7532 31892 7588 31902
rect 7420 31836 7532 31892
rect 7420 31220 7476 31836
rect 7532 31826 7588 31836
rect 7868 31890 7924 34300
rect 7980 33460 8036 33470
rect 7980 33366 8036 33404
rect 7868 31838 7870 31890
rect 7922 31838 7924 31890
rect 7868 31826 7924 31838
rect 8092 33122 8148 34412
rect 8988 34132 9044 34142
rect 8988 34038 9044 34076
rect 8876 33906 8932 33918
rect 8876 33854 8878 33906
rect 8930 33854 8932 33906
rect 8876 33572 8932 33854
rect 8316 33348 8372 33358
rect 8876 33348 8932 33516
rect 8316 33346 8932 33348
rect 8316 33294 8318 33346
rect 8370 33294 8932 33346
rect 8316 33292 8932 33294
rect 8988 33796 9044 33806
rect 8316 33282 8372 33292
rect 8988 33236 9044 33740
rect 8092 33070 8094 33122
rect 8146 33070 8148 33122
rect 7980 31780 8036 31790
rect 8092 31780 8148 33070
rect 8764 33180 9044 33236
rect 8764 32562 8820 33180
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 32498 8820 32510
rect 9212 33122 9268 33134
rect 9212 33070 9214 33122
rect 9266 33070 9268 33122
rect 7980 31778 8148 31780
rect 7980 31726 7982 31778
rect 8034 31726 8148 31778
rect 7980 31724 8148 31726
rect 7980 31714 8036 31724
rect 7532 31556 7588 31566
rect 7532 31554 7700 31556
rect 7532 31502 7534 31554
rect 7586 31502 7700 31554
rect 7532 31500 7700 31502
rect 7532 31490 7588 31500
rect 7532 31220 7588 31230
rect 7420 31218 7588 31220
rect 7420 31166 7534 31218
rect 7586 31166 7588 31218
rect 7420 31164 7588 31166
rect 7196 30994 7476 30996
rect 7196 30942 7198 30994
rect 7250 30942 7476 30994
rect 7196 30940 7476 30942
rect 7196 30930 7252 30940
rect 7308 30770 7364 30782
rect 7308 30718 7310 30770
rect 7362 30718 7364 30770
rect 7196 30324 7252 30334
rect 7308 30324 7364 30718
rect 7252 30268 7364 30324
rect 7196 30230 7252 30268
rect 7140 29708 7252 29764
rect 7084 29698 7140 29708
rect 6412 29202 6692 29204
rect 6412 29150 6638 29202
rect 6690 29150 6692 29202
rect 6412 29148 6692 29150
rect 6412 28866 6468 29148
rect 6636 29138 6692 29148
rect 6748 29148 7028 29204
rect 6412 28814 6414 28866
rect 6466 28814 6468 28866
rect 6412 28802 6468 28814
rect 6412 28532 6468 28542
rect 6188 28084 6244 28094
rect 6188 27990 6244 28028
rect 5852 27860 5908 27870
rect 5852 27858 6020 27860
rect 5852 27806 5854 27858
rect 5906 27806 6020 27858
rect 5852 27804 6020 27806
rect 5852 27794 5908 27804
rect 5964 27412 6020 27804
rect 5628 27356 5796 27412
rect 5292 27122 5348 27132
rect 5180 26852 5572 26908
rect 5068 24894 5070 24946
rect 5122 24894 5124 24946
rect 5068 24882 5124 24894
rect 5404 25508 5460 25518
rect 4620 24724 4676 24734
rect 4620 24610 4676 24668
rect 5404 24724 5460 25452
rect 5404 24630 5460 24668
rect 4620 24558 4622 24610
rect 4674 24558 4676 24610
rect 4620 24546 4676 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 2940 24110 2942 24162
rect 2994 24110 2996 24162
rect 2940 24098 2996 24110
rect 5516 23828 5572 26852
rect 5740 26402 5796 27356
rect 5740 26350 5742 26402
rect 5794 26350 5796 26402
rect 5628 25508 5684 25518
rect 5628 25414 5684 25452
rect 5740 24948 5796 26350
rect 5852 27356 6020 27412
rect 5852 26516 5908 27356
rect 6076 27300 6132 27916
rect 5964 27244 6132 27300
rect 5964 26908 6020 27244
rect 5964 26852 6132 26908
rect 5852 25506 5908 26460
rect 6076 26402 6132 26852
rect 6076 26350 6078 26402
rect 6130 26350 6132 26402
rect 6076 26292 6132 26350
rect 6076 26226 6132 26236
rect 6412 25844 6468 28476
rect 6636 28084 6692 28094
rect 6636 27970 6692 28028
rect 6636 27918 6638 27970
rect 6690 27918 6692 27970
rect 6636 27906 6692 27918
rect 6524 27858 6580 27870
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 27636 6580 27806
rect 6524 27570 6580 27580
rect 6636 27300 6692 27310
rect 6636 27206 6692 27244
rect 6524 27188 6580 27198
rect 6524 27094 6580 27132
rect 6636 26516 6692 26526
rect 6636 26422 6692 26460
rect 6524 26292 6580 26302
rect 6524 26198 6580 26236
rect 6748 26292 6804 29148
rect 7196 28532 7252 29708
rect 7196 28466 7252 28476
rect 7308 27970 7364 27982
rect 7308 27918 7310 27970
rect 7362 27918 7364 27970
rect 6972 27860 7028 27870
rect 7196 27860 7252 27870
rect 6972 27858 7252 27860
rect 6972 27806 6974 27858
rect 7026 27806 7198 27858
rect 7250 27806 7252 27858
rect 6972 27804 7252 27806
rect 6972 27794 7028 27804
rect 7196 27794 7252 27804
rect 6860 27748 6916 27758
rect 6860 27654 6916 27692
rect 7308 27300 7364 27918
rect 7308 27234 7364 27244
rect 7420 26908 7476 30940
rect 7532 30770 7588 31164
rect 7532 30718 7534 30770
rect 7586 30718 7588 30770
rect 7532 30706 7588 30718
rect 7532 28084 7588 28094
rect 7532 27990 7588 28028
rect 7196 26852 7476 26908
rect 7644 26908 7700 31500
rect 7756 31554 7812 31566
rect 7756 31502 7758 31554
rect 7810 31502 7812 31554
rect 7756 30212 7812 31502
rect 7756 30146 7812 30156
rect 8204 31556 8260 31566
rect 8204 28642 8260 31500
rect 8204 28590 8206 28642
rect 8258 28590 8260 28642
rect 8204 28578 8260 28590
rect 8316 30324 8372 30334
rect 8316 28082 8372 30268
rect 8652 30212 8708 30222
rect 8428 30100 8484 30110
rect 8428 28644 8484 30044
rect 8652 29538 8708 30156
rect 8652 29486 8654 29538
rect 8706 29486 8708 29538
rect 8652 29474 8708 29486
rect 8876 29538 8932 29550
rect 8876 29486 8878 29538
rect 8930 29486 8932 29538
rect 8876 29428 8932 29486
rect 8876 29362 8932 29372
rect 8988 29316 9044 29326
rect 8988 29222 9044 29260
rect 8428 28550 8484 28588
rect 8540 28642 8596 28654
rect 8540 28590 8542 28642
rect 8594 28590 8596 28642
rect 8316 28030 8318 28082
rect 8370 28030 8372 28082
rect 7756 27972 7812 27982
rect 7756 27878 7812 27916
rect 8316 27636 8372 28030
rect 8540 27860 8596 28590
rect 8540 27794 8596 27804
rect 8988 28418 9044 28430
rect 8988 28366 8990 28418
rect 9042 28366 9044 28418
rect 8316 27570 8372 27580
rect 7644 26852 7924 26908
rect 6972 26292 7028 26302
rect 6748 26290 6916 26292
rect 6748 26238 6750 26290
rect 6802 26238 6916 26290
rect 6748 26236 6916 26238
rect 6748 26226 6804 26236
rect 6412 25788 6804 25844
rect 5852 25454 5854 25506
rect 5906 25454 5908 25506
rect 5852 25442 5908 25454
rect 6076 25620 6132 25630
rect 6636 25620 6692 25630
rect 6076 25506 6132 25564
rect 6076 25454 6078 25506
rect 6130 25454 6132 25506
rect 5964 25284 6020 25294
rect 5964 25190 6020 25228
rect 5964 24948 6020 24958
rect 5740 24946 6020 24948
rect 5740 24894 5966 24946
rect 6018 24894 6020 24946
rect 5740 24892 6020 24894
rect 5964 24882 6020 24892
rect 5628 24724 5684 24734
rect 6076 24724 6132 25454
rect 6300 25618 6692 25620
rect 6300 25566 6638 25618
rect 6690 25566 6692 25618
rect 6300 25564 6692 25566
rect 6300 25506 6356 25564
rect 6636 25554 6692 25564
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 6300 25442 6356 25454
rect 6748 25396 6804 25788
rect 5628 24722 6132 24724
rect 5628 24670 5630 24722
rect 5682 24670 6132 24722
rect 5628 24668 6132 24670
rect 6412 25394 6804 25396
rect 6412 25342 6750 25394
rect 6802 25342 6804 25394
rect 6412 25340 6804 25342
rect 5628 24658 5684 24668
rect 5628 23828 5684 23838
rect 4844 23826 5684 23828
rect 4844 23774 5630 23826
rect 5682 23774 5684 23826
rect 4844 23772 5684 23774
rect 2716 23716 2772 23726
rect 2716 23622 2772 23660
rect 3388 23716 3444 23726
rect 3500 23716 3556 23726
rect 3444 23714 3556 23716
rect 3444 23662 3502 23714
rect 3554 23662 3556 23714
rect 3444 23660 3556 23662
rect 1708 22318 1710 22370
rect 1762 22318 1764 22370
rect 1708 20244 1764 22318
rect 2492 22260 2548 22270
rect 2492 22258 2660 22260
rect 2492 22206 2494 22258
rect 2546 22206 2660 22258
rect 2492 22204 2660 22206
rect 2492 22194 2548 22204
rect 2604 21474 2660 22204
rect 2940 22148 2996 22158
rect 2604 21422 2606 21474
rect 2658 21422 2660 21474
rect 2604 21410 2660 21422
rect 2716 21698 2772 21710
rect 2716 21646 2718 21698
rect 2770 21646 2772 21698
rect 1708 19234 1764 20188
rect 2716 20132 2772 21646
rect 2940 21698 2996 22092
rect 2940 21646 2942 21698
rect 2994 21646 2996 21698
rect 2940 21634 2996 21646
rect 3388 21476 3444 23660
rect 3500 23650 3556 23660
rect 4844 23266 4900 23772
rect 5628 23762 5684 23772
rect 5964 23716 6020 23726
rect 4844 23214 4846 23266
rect 4898 23214 4900 23266
rect 4844 23202 4900 23214
rect 5068 23266 5124 23278
rect 5068 23214 5070 23266
rect 5122 23214 5124 23266
rect 4620 23042 4676 23054
rect 4620 22990 4622 23042
rect 4674 22990 4676 23042
rect 4620 22932 4676 22990
rect 4620 22876 4900 22932
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4620 22484 4676 22494
rect 4844 22484 4900 22876
rect 5068 22484 5124 23214
rect 5964 23156 6020 23660
rect 6412 23378 6468 25340
rect 6748 25330 6804 25340
rect 6860 24948 6916 26236
rect 6972 25730 7028 26236
rect 6972 25678 6974 25730
rect 7026 25678 7028 25730
rect 6972 25666 7028 25678
rect 7196 26290 7252 26852
rect 7196 26238 7198 26290
rect 7250 26238 7252 26290
rect 6972 24948 7028 24958
rect 6860 24946 7028 24948
rect 6860 24894 6974 24946
rect 7026 24894 7028 24946
rect 6860 24892 7028 24894
rect 6972 24882 7028 24892
rect 6636 24722 6692 24734
rect 6636 24670 6638 24722
rect 6690 24670 6692 24722
rect 6636 23716 6692 24670
rect 6636 23650 6692 23660
rect 7196 23492 7252 26238
rect 7196 23426 7252 23436
rect 7868 23938 7924 26852
rect 8988 25506 9044 28366
rect 9212 26908 9268 33070
rect 9324 30210 9380 34860
rect 9884 34850 9940 34860
rect 9660 34692 9716 34702
rect 9548 34636 9660 34692
rect 9548 33796 9604 34636
rect 9660 34626 9716 34636
rect 9996 34356 10052 35534
rect 10220 35026 10276 36318
rect 10668 36260 10724 36270
rect 10668 35476 10724 36204
rect 10668 35410 10724 35420
rect 10220 34974 10222 35026
rect 10274 34974 10276 35026
rect 10220 34962 10276 34974
rect 10332 34916 10388 34926
rect 9884 34300 10052 34356
rect 10108 34690 10164 34702
rect 10108 34638 10110 34690
rect 10162 34638 10164 34690
rect 9660 33908 9716 33946
rect 9660 33842 9716 33852
rect 9772 33906 9828 33918
rect 9772 33854 9774 33906
rect 9826 33854 9828 33906
rect 9548 32788 9604 33740
rect 9660 33684 9716 33694
rect 9660 33124 9716 33628
rect 9772 33572 9828 33854
rect 9884 33684 9940 34300
rect 10108 34242 10164 34638
rect 10108 34190 10110 34242
rect 10162 34190 10164 34242
rect 10108 34178 10164 34190
rect 9996 34020 10052 34030
rect 10332 34020 10388 34860
rect 10444 34690 10500 34702
rect 10444 34638 10446 34690
rect 10498 34638 10500 34690
rect 10444 34356 10500 34638
rect 11004 34692 11060 34702
rect 11004 34598 11060 34636
rect 10444 34290 10500 34300
rect 9996 34018 10388 34020
rect 9996 33966 9998 34018
rect 10050 33966 10388 34018
rect 9996 33964 10388 33966
rect 10892 34018 10948 34030
rect 10892 33966 10894 34018
rect 10946 33966 10948 34018
rect 9996 33954 10052 33964
rect 9884 33628 10052 33684
rect 9772 33348 9828 33516
rect 9996 33458 10052 33628
rect 9996 33406 9998 33458
rect 10050 33406 10052 33458
rect 9996 33394 10052 33406
rect 9884 33348 9940 33358
rect 9772 33346 9940 33348
rect 9772 33294 9886 33346
rect 9938 33294 9940 33346
rect 9772 33292 9940 33294
rect 9884 33282 9940 33292
rect 10220 33346 10276 33358
rect 10220 33294 10222 33346
rect 10274 33294 10276 33346
rect 10220 33124 10276 33294
rect 9660 33068 9940 33124
rect 9660 32788 9716 32798
rect 9548 32786 9716 32788
rect 9548 32734 9662 32786
rect 9714 32734 9716 32786
rect 9548 32732 9716 32734
rect 9660 32722 9716 32732
rect 9436 32452 9492 32462
rect 9436 31892 9492 32396
rect 9436 31890 9828 31892
rect 9436 31838 9438 31890
rect 9490 31838 9828 31890
rect 9436 31836 9828 31838
rect 9436 31826 9492 31836
rect 9772 31778 9828 31836
rect 9772 31726 9774 31778
rect 9826 31726 9828 31778
rect 9772 31714 9828 31726
rect 9884 31556 9940 33068
rect 10220 33058 10276 33068
rect 10892 31892 10948 33966
rect 11004 33346 11060 33358
rect 11004 33294 11006 33346
rect 11058 33294 11060 33346
rect 11004 33124 11060 33294
rect 11004 33058 11060 33068
rect 10892 31826 10948 31836
rect 10556 31668 10612 31678
rect 9772 31500 9940 31556
rect 10108 31666 10612 31668
rect 10108 31614 10558 31666
rect 10610 31614 10612 31666
rect 10108 31612 10612 31614
rect 9772 30994 9828 31500
rect 10108 31218 10164 31612
rect 10556 31602 10612 31612
rect 10108 31166 10110 31218
rect 10162 31166 10164 31218
rect 10108 31154 10164 31166
rect 9772 30942 9774 30994
rect 9826 30942 9828 30994
rect 9772 30930 9828 30942
rect 9884 30996 9940 31006
rect 9884 30434 9940 30940
rect 9884 30382 9886 30434
rect 9938 30382 9940 30434
rect 9884 30370 9940 30382
rect 9996 30994 10052 31006
rect 9996 30942 9998 30994
rect 10050 30942 10052 30994
rect 9324 30158 9326 30210
rect 9378 30158 9380 30210
rect 9324 28084 9380 30158
rect 9548 29986 9604 29998
rect 9548 29934 9550 29986
rect 9602 29934 9604 29986
rect 9548 29428 9604 29934
rect 9772 29986 9828 29998
rect 9772 29934 9774 29986
rect 9826 29934 9828 29986
rect 9548 29362 9604 29372
rect 9660 29538 9716 29550
rect 9660 29486 9662 29538
rect 9714 29486 9716 29538
rect 9660 28756 9716 29486
rect 9772 28868 9828 29934
rect 9996 29650 10052 30942
rect 10220 30996 10276 31006
rect 10220 30902 10276 30940
rect 9996 29598 9998 29650
rect 10050 29598 10052 29650
rect 9996 29586 10052 29598
rect 10108 29652 10164 29662
rect 10108 29650 11060 29652
rect 10108 29598 10110 29650
rect 10162 29598 11060 29650
rect 10108 29596 11060 29598
rect 10108 29586 10164 29596
rect 9884 29426 9940 29438
rect 9884 29374 9886 29426
rect 9938 29374 9940 29426
rect 9884 29316 9940 29374
rect 9884 29250 9940 29260
rect 10444 29426 10500 29438
rect 10444 29374 10446 29426
rect 10498 29374 10500 29426
rect 10444 29316 10500 29374
rect 10444 29250 10500 29260
rect 10780 29428 10836 29438
rect 10108 28868 10164 28878
rect 9772 28866 10164 28868
rect 9772 28814 10110 28866
rect 10162 28814 10164 28866
rect 9772 28812 10164 28814
rect 10108 28802 10164 28812
rect 9660 28690 9716 28700
rect 10220 28756 10276 28766
rect 10220 28662 10276 28700
rect 10668 28532 10724 28542
rect 9380 28028 9604 28084
rect 9324 28018 9380 28028
rect 9212 26852 9380 26908
rect 9324 25620 9380 26852
rect 9548 26514 9604 28028
rect 10332 27970 10388 27982
rect 10332 27918 10334 27970
rect 10386 27918 10388 27970
rect 10332 27076 10388 27918
rect 10668 27970 10724 28476
rect 10668 27918 10670 27970
rect 10722 27918 10724 27970
rect 10668 27906 10724 27918
rect 10780 27076 10836 29372
rect 11004 29426 11060 29596
rect 11004 29374 11006 29426
rect 11058 29374 11060 29426
rect 10892 29316 10948 29326
rect 10892 29222 10948 29260
rect 11004 27300 11060 29374
rect 11004 27234 11060 27244
rect 11004 27076 11060 27086
rect 10332 27074 11060 27076
rect 10332 27022 11006 27074
rect 11058 27022 11060 27074
rect 10332 27020 11060 27022
rect 11004 27010 11060 27020
rect 9548 26462 9550 26514
rect 9602 26462 9604 26514
rect 9548 26450 9604 26462
rect 11004 26852 11060 26862
rect 9772 26290 9828 26302
rect 9772 26238 9774 26290
rect 9826 26238 9828 26290
rect 9772 25956 9828 26238
rect 11004 26068 11060 26796
rect 11004 26002 11060 26012
rect 9324 25554 9380 25564
rect 9548 25900 9828 25956
rect 8988 25454 8990 25506
rect 9042 25454 9044 25506
rect 8988 25442 9044 25454
rect 9436 25508 9492 25518
rect 9436 25394 9492 25452
rect 9436 25342 9438 25394
rect 9490 25342 9492 25394
rect 9436 25330 9492 25342
rect 9548 25396 9604 25900
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 6412 23326 6414 23378
rect 6466 23326 6468 23378
rect 6188 23156 6244 23166
rect 5964 23154 6244 23156
rect 5964 23102 6190 23154
rect 6242 23102 6244 23154
rect 5964 23100 6244 23102
rect 5180 22932 5236 22942
rect 5180 22930 5348 22932
rect 5180 22878 5182 22930
rect 5234 22878 5348 22930
rect 5180 22876 5348 22878
rect 5180 22866 5236 22876
rect 4620 22482 5124 22484
rect 4620 22430 4622 22482
rect 4674 22430 5070 22482
rect 5122 22430 5124 22482
rect 4620 22428 5124 22430
rect 4620 22418 4676 22428
rect 5068 22372 5124 22428
rect 5180 22372 5236 22382
rect 5068 22316 5180 22372
rect 5180 22306 5236 22316
rect 5292 22036 5348 22876
rect 6188 22484 6244 23100
rect 5292 21970 5348 21980
rect 5628 22428 6244 22484
rect 5404 21812 5460 21822
rect 5404 21718 5460 21756
rect 5628 21588 5684 22428
rect 5852 22260 5908 22270
rect 6300 22260 6356 22270
rect 5852 22166 5908 22204
rect 6188 22258 6356 22260
rect 6188 22206 6302 22258
rect 6354 22206 6356 22258
rect 6188 22204 6356 22206
rect 5516 21586 5684 21588
rect 5516 21534 5630 21586
rect 5682 21534 5684 21586
rect 5516 21532 5684 21534
rect 3388 21474 3556 21476
rect 3388 21422 3390 21474
rect 3442 21422 3556 21474
rect 3388 21420 3556 21422
rect 3388 21410 3444 21420
rect 3052 20580 3108 20590
rect 2828 20132 2884 20142
rect 2716 20076 2828 20132
rect 2828 20038 2884 20076
rect 3052 20130 3108 20524
rect 3052 20078 3054 20130
rect 3106 20078 3108 20130
rect 3052 20066 3108 20078
rect 3500 20132 3556 21420
rect 4844 21474 4900 21486
rect 4844 21422 4846 21474
rect 4898 21422 4900 21474
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 20244 4900 21422
rect 4900 20188 5124 20244
rect 4844 20178 4900 20188
rect 3500 20038 3556 20076
rect 4956 20020 5012 20030
rect 2716 19796 2772 19806
rect 2492 19794 2772 19796
rect 2492 19742 2718 19794
rect 2770 19742 2772 19794
rect 2492 19740 2772 19742
rect 2492 19346 2548 19740
rect 2716 19730 2772 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2492 19282 2548 19294
rect 4620 19348 4676 19358
rect 4956 19348 5012 19964
rect 4620 19346 5012 19348
rect 4620 19294 4622 19346
rect 4674 19294 5012 19346
rect 4620 19292 5012 19294
rect 5068 19348 5124 20188
rect 5180 20020 5236 20030
rect 5180 19926 5236 19964
rect 5180 19348 5236 19358
rect 5068 19346 5236 19348
rect 5068 19294 5182 19346
rect 5234 19294 5236 19346
rect 5068 19292 5236 19294
rect 4620 19282 4676 19292
rect 5180 19282 5236 19292
rect 1708 19182 1710 19234
rect 1762 19182 1764 19234
rect 1708 19170 1764 19182
rect 5516 18564 5572 21532
rect 5628 21522 5684 21532
rect 5740 22146 5796 22158
rect 5740 22094 5742 22146
rect 5794 22094 5796 22146
rect 5740 21810 5796 22094
rect 5964 22148 6020 22158
rect 5964 22054 6020 22092
rect 6076 22146 6132 22158
rect 6076 22094 6078 22146
rect 6130 22094 6132 22146
rect 6076 22036 6132 22094
rect 6076 21970 6132 21980
rect 5740 21758 5742 21810
rect 5794 21758 5796 21810
rect 5628 20804 5684 20814
rect 5740 20804 5796 21758
rect 5852 21700 5908 21710
rect 5852 21606 5908 21644
rect 6188 21700 6244 22204
rect 6300 22194 6356 22204
rect 6188 21634 6244 21644
rect 6412 21588 6468 23326
rect 7532 23044 7588 23054
rect 7084 22484 7140 22494
rect 7532 22484 7588 22988
rect 7084 22482 7588 22484
rect 7084 22430 7086 22482
rect 7138 22430 7588 22482
rect 7084 22428 7588 22430
rect 7084 22372 7140 22428
rect 7084 22306 7140 22316
rect 7420 22260 7476 22270
rect 7196 22258 7476 22260
rect 7196 22206 7422 22258
rect 7474 22206 7476 22258
rect 7196 22204 7476 22206
rect 6524 21588 6580 21598
rect 6412 21586 6580 21588
rect 6412 21534 6526 21586
rect 6578 21534 6580 21586
rect 6412 21532 6580 21534
rect 6524 21522 6580 21532
rect 6636 21588 6692 21598
rect 7084 21588 7140 21598
rect 6636 21494 6692 21532
rect 6748 21586 7140 21588
rect 6748 21534 7086 21586
rect 7138 21534 7140 21586
rect 6748 21532 7140 21534
rect 6300 21476 6356 21486
rect 6356 21420 6468 21476
rect 6300 21382 6356 21420
rect 5628 20802 5796 20804
rect 5628 20750 5630 20802
rect 5682 20750 5796 20802
rect 5628 20748 5796 20750
rect 6188 21362 6244 21374
rect 6188 21310 6190 21362
rect 6242 21310 6244 21362
rect 6188 20802 6244 21310
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 5628 20738 5684 20748
rect 6188 20738 6244 20750
rect 6412 20916 6468 21420
rect 6636 21028 6692 21038
rect 6748 21028 6804 21532
rect 7084 21522 7140 21532
rect 7196 21476 7252 22204
rect 7420 22194 7476 22204
rect 7532 22258 7588 22428
rect 7532 22206 7534 22258
rect 7586 22206 7588 22258
rect 7532 22194 7588 22206
rect 7644 22372 7700 22382
rect 7308 21700 7364 21710
rect 7308 21606 7364 21644
rect 7420 21700 7476 21710
rect 7644 21700 7700 22316
rect 7756 22260 7812 22270
rect 7756 22166 7812 22204
rect 7420 21698 7700 21700
rect 7420 21646 7422 21698
rect 7474 21646 7700 21698
rect 7420 21644 7700 21646
rect 7868 21812 7924 23886
rect 8988 25282 9044 25294
rect 8988 25230 8990 25282
rect 9042 25230 9044 25282
rect 8092 23714 8148 23726
rect 8092 23662 8094 23714
rect 8146 23662 8148 23714
rect 8092 23492 8148 23662
rect 8092 23426 8148 23436
rect 8316 22596 8372 22606
rect 8316 22502 8372 22540
rect 8988 22594 9044 25230
rect 9548 22708 9604 25340
rect 9660 25620 9716 25630
rect 9660 25394 9716 25564
rect 9660 25342 9662 25394
rect 9714 25342 9716 25394
rect 9660 25330 9716 25342
rect 10332 25396 10388 25406
rect 10332 25302 10388 25340
rect 10668 25396 10724 25406
rect 10668 25302 10724 25340
rect 11116 25284 11172 38780
rect 11564 38668 11620 39452
rect 11676 39394 11732 39406
rect 11676 39342 11678 39394
rect 11730 39342 11732 39394
rect 11676 39060 11732 39342
rect 11676 38994 11732 39004
rect 11564 38612 11732 38668
rect 11564 35028 11620 35038
rect 11676 35028 11732 38612
rect 11788 36932 11844 43484
rect 12012 42084 12068 43820
rect 12124 44098 12180 44110
rect 12124 44046 12126 44098
rect 12178 44046 12180 44098
rect 12124 43708 12180 44046
rect 12124 43652 12516 43708
rect 12460 42756 12516 43652
rect 12348 42754 12516 42756
rect 12348 42702 12462 42754
rect 12514 42702 12516 42754
rect 12348 42700 12516 42702
rect 12236 42084 12292 42094
rect 12012 42028 12236 42084
rect 12236 42018 12292 42028
rect 12348 41970 12404 42700
rect 12460 42690 12516 42700
rect 12348 41918 12350 41970
rect 12402 41918 12404 41970
rect 12124 41858 12180 41870
rect 12124 41806 12126 41858
rect 12178 41806 12180 41858
rect 12124 41076 12180 41806
rect 12348 41186 12404 41918
rect 12348 41134 12350 41186
rect 12402 41134 12404 41186
rect 12348 41122 12404 41134
rect 12572 42530 12628 42542
rect 12572 42478 12574 42530
rect 12626 42478 12628 42530
rect 12124 41010 12180 41020
rect 12572 41076 12628 42478
rect 12796 42532 12852 42542
rect 12796 42530 13412 42532
rect 12796 42478 12798 42530
rect 12850 42478 13412 42530
rect 12796 42476 13412 42478
rect 12796 42466 12852 42476
rect 12684 42252 13188 42308
rect 12684 42194 12740 42252
rect 12684 42142 12686 42194
rect 12738 42142 12740 42194
rect 12684 42130 12740 42142
rect 13132 42196 13188 42252
rect 13244 42196 13300 42206
rect 13132 42194 13300 42196
rect 13132 42142 13246 42194
rect 13298 42142 13300 42194
rect 13132 42140 13300 42142
rect 13244 42130 13300 42140
rect 13020 42084 13076 42094
rect 13020 41990 13076 42028
rect 12908 41972 12964 41982
rect 13356 41972 13412 42476
rect 13468 41972 13524 41982
rect 13356 41970 13524 41972
rect 13356 41918 13470 41970
rect 13522 41918 13524 41970
rect 13356 41916 13524 41918
rect 12908 41878 12964 41916
rect 12684 41188 12740 41198
rect 12684 41094 12740 41132
rect 13468 41186 13524 41916
rect 13468 41134 13470 41186
rect 13522 41134 13524 41186
rect 13468 41122 13524 41134
rect 12572 41010 12628 41020
rect 12908 41076 12964 41086
rect 12908 40982 12964 41020
rect 13020 40964 13076 40974
rect 13020 40962 13300 40964
rect 13020 40910 13022 40962
rect 13074 40910 13300 40962
rect 13020 40908 13300 40910
rect 13020 40898 13076 40908
rect 11788 36866 11844 36876
rect 11900 40404 11956 40414
rect 11788 35924 11844 35934
rect 11788 35698 11844 35868
rect 11788 35646 11790 35698
rect 11842 35646 11844 35698
rect 11788 35634 11844 35646
rect 11340 35026 11732 35028
rect 11340 34974 11566 35026
rect 11618 34974 11732 35026
rect 11340 34972 11732 34974
rect 11340 34354 11396 34972
rect 11564 34962 11620 34972
rect 11900 34468 11956 40348
rect 13244 39508 13300 40908
rect 13468 39508 13524 39518
rect 13244 39506 13524 39508
rect 13244 39454 13470 39506
rect 13522 39454 13524 39506
rect 13244 39452 13524 39454
rect 13580 39508 13636 44156
rect 13692 41972 13748 41982
rect 13692 41188 13748 41916
rect 13692 41094 13748 41132
rect 13804 39844 13860 48972
rect 16268 47460 16324 47470
rect 16268 47366 16324 47404
rect 17948 47460 18004 50540
rect 19628 50036 19684 50652
rect 19740 50642 19796 50652
rect 23100 50708 23156 50718
rect 23100 50614 23156 50652
rect 26124 50708 26180 50718
rect 20188 50596 20244 50606
rect 21196 50596 21252 50606
rect 20188 50502 20244 50540
rect 20524 50594 21252 50596
rect 20524 50542 21198 50594
rect 21250 50542 21252 50594
rect 20524 50540 21252 50542
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19628 49810 19684 49980
rect 20412 50036 20468 50046
rect 19628 49758 19630 49810
rect 19682 49758 19684 49810
rect 19628 49746 19684 49758
rect 19852 49924 19908 49934
rect 19852 49810 19908 49868
rect 19852 49758 19854 49810
rect 19906 49758 19908 49810
rect 19852 49746 19908 49758
rect 20076 49588 20132 49598
rect 20076 49494 20132 49532
rect 20412 48914 20468 49980
rect 20524 50034 20580 50540
rect 21196 50530 21252 50540
rect 21532 50594 21588 50606
rect 21532 50542 21534 50594
rect 21586 50542 21588 50594
rect 21420 50484 21476 50494
rect 21420 50390 21476 50428
rect 20524 49982 20526 50034
rect 20578 49982 20580 50034
rect 20524 49970 20580 49982
rect 21196 50036 21252 50046
rect 21196 49942 21252 49980
rect 21308 49812 21364 49822
rect 21308 49718 21364 49756
rect 21196 49588 21252 49598
rect 21532 49588 21588 50542
rect 24332 50594 24388 50606
rect 24332 50542 24334 50594
rect 24386 50542 24388 50594
rect 21868 50484 21924 50494
rect 21868 50390 21924 50428
rect 22092 50484 22148 50494
rect 22092 50148 22148 50428
rect 22988 50484 23044 50494
rect 22988 50390 23044 50428
rect 23212 50482 23268 50494
rect 23212 50430 23214 50482
rect 23266 50430 23268 50482
rect 22764 50372 22820 50382
rect 22764 50370 22932 50372
rect 22764 50318 22766 50370
rect 22818 50318 22932 50370
rect 22764 50316 22932 50318
rect 22764 50306 22820 50316
rect 21868 50092 22148 50148
rect 21868 50034 21924 50092
rect 21868 49982 21870 50034
rect 21922 49982 21924 50034
rect 21868 49970 21924 49982
rect 21980 49922 22036 49934
rect 21980 49870 21982 49922
rect 22034 49870 22036 49922
rect 21980 49700 22036 49870
rect 21868 49644 22036 49700
rect 21196 49586 21588 49588
rect 21196 49534 21198 49586
rect 21250 49534 21588 49586
rect 21196 49532 21588 49534
rect 21644 49588 21700 49598
rect 21756 49588 21812 49598
rect 21700 49586 21812 49588
rect 21700 49534 21758 49586
rect 21810 49534 21812 49586
rect 21700 49532 21812 49534
rect 21196 49522 21252 49532
rect 20748 49028 20804 49038
rect 20748 48934 20804 48972
rect 21644 49026 21700 49532
rect 21756 49522 21812 49532
rect 21644 48974 21646 49026
rect 21698 48974 21700 49026
rect 20412 48862 20414 48914
rect 20466 48862 20468 48914
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 16940 47348 16996 47358
rect 16940 47254 16996 47292
rect 17948 46900 18004 47404
rect 19068 47570 19124 47582
rect 19068 47518 19070 47570
rect 19122 47518 19124 47570
rect 19068 47236 19124 47518
rect 20300 47346 20356 47358
rect 20300 47294 20302 47346
rect 20354 47294 20356 47346
rect 19404 47236 19460 47246
rect 19740 47236 19796 47246
rect 19068 47234 19460 47236
rect 19068 47182 19406 47234
rect 19458 47182 19460 47234
rect 19068 47180 19460 47182
rect 19292 46900 19348 46910
rect 18004 46844 18116 46900
rect 17948 46806 18004 46844
rect 15820 46676 15876 46686
rect 15820 46562 15876 46620
rect 15820 46510 15822 46562
rect 15874 46510 15876 46562
rect 13916 45780 13972 45790
rect 13916 45106 13972 45724
rect 14812 45780 14868 45790
rect 14812 45330 14868 45724
rect 14812 45278 14814 45330
rect 14866 45278 14868 45330
rect 14812 45266 14868 45278
rect 13916 45054 13918 45106
rect 13970 45054 13972 45106
rect 13916 45042 13972 45054
rect 14252 45108 14308 45118
rect 14252 45014 14308 45052
rect 14364 44994 14420 45006
rect 14364 44942 14366 44994
rect 14418 44942 14420 44994
rect 14140 44212 14196 44222
rect 14364 44212 14420 44942
rect 14196 44156 14420 44212
rect 14476 44322 14532 44334
rect 14476 44270 14478 44322
rect 14530 44270 14532 44322
rect 14476 44212 14532 44270
rect 14140 44146 14196 44156
rect 14476 44146 14532 44156
rect 15148 44212 15204 44222
rect 14700 44098 14756 44110
rect 14700 44046 14702 44098
rect 14754 44046 14756 44098
rect 14700 43988 14756 44046
rect 14700 43922 14756 43932
rect 15148 44098 15204 44156
rect 15148 44046 15150 44098
rect 15202 44046 15204 44098
rect 15148 43708 15204 44046
rect 14924 43652 15204 43708
rect 14812 42754 14868 42766
rect 14812 42702 14814 42754
rect 14866 42702 14868 42754
rect 14812 42532 14868 42702
rect 14812 42466 14868 42476
rect 14028 41412 14084 41422
rect 14028 41410 14196 41412
rect 14028 41358 14030 41410
rect 14082 41358 14196 41410
rect 14028 41356 14196 41358
rect 14028 41346 14084 41356
rect 14140 41300 14196 41356
rect 14812 41300 14868 41310
rect 14924 41300 14980 43652
rect 15484 43316 15540 43326
rect 15484 42866 15540 43260
rect 15484 42814 15486 42866
rect 15538 42814 15540 42866
rect 15484 42802 15540 42814
rect 14140 41298 14980 41300
rect 14140 41246 14814 41298
rect 14866 41246 14980 41298
rect 14140 41244 14980 41246
rect 14812 41234 14868 41244
rect 14028 41188 14084 41198
rect 14028 41186 14532 41188
rect 14028 41134 14030 41186
rect 14082 41134 14532 41186
rect 14028 41132 14532 41134
rect 13804 39778 13860 39788
rect 13916 40962 13972 40974
rect 13916 40910 13918 40962
rect 13970 40910 13972 40962
rect 13916 39842 13972 40910
rect 13916 39790 13918 39842
rect 13970 39790 13972 39842
rect 13916 39778 13972 39790
rect 13804 39620 13860 39630
rect 14028 39620 14084 41132
rect 14252 40178 14308 40190
rect 14252 40126 14254 40178
rect 14306 40126 14308 40178
rect 13804 39618 14084 39620
rect 13804 39566 13806 39618
rect 13858 39566 14084 39618
rect 13804 39564 14084 39566
rect 14140 39844 14196 39854
rect 13804 39554 13860 39564
rect 13580 39452 13748 39508
rect 13468 39442 13524 39452
rect 12124 39396 12180 39406
rect 12012 39284 12068 39294
rect 12012 35476 12068 39228
rect 12124 38834 12180 39340
rect 12796 38948 12852 38958
rect 12796 38854 12852 38892
rect 12124 38782 12126 38834
rect 12178 38782 12180 38834
rect 12124 38770 12180 38782
rect 13692 37266 13748 39452
rect 13916 39394 13972 39406
rect 13916 39342 13918 39394
rect 13970 39342 13972 39394
rect 13916 38948 13972 39342
rect 13916 38882 13972 38892
rect 14140 38724 14196 39788
rect 13692 37214 13694 37266
rect 13746 37214 13748 37266
rect 13692 37202 13748 37214
rect 13916 38668 14196 38724
rect 14252 39618 14308 40126
rect 14476 39844 14532 41132
rect 14588 40290 14644 40302
rect 14588 40238 14590 40290
rect 14642 40238 14644 40290
rect 14588 40178 14644 40238
rect 14588 40126 14590 40178
rect 14642 40126 14644 40178
rect 14588 40114 14644 40126
rect 14588 39844 14644 39854
rect 14476 39842 14644 39844
rect 14476 39790 14590 39842
rect 14642 39790 14644 39842
rect 14476 39788 14644 39790
rect 14588 39778 14644 39788
rect 14252 39566 14254 39618
rect 14306 39566 14308 39618
rect 14252 38668 14308 39566
rect 15484 39732 15540 39742
rect 15484 39618 15540 39676
rect 15484 39566 15486 39618
rect 15538 39566 15540 39618
rect 14700 39506 14756 39518
rect 14700 39454 14702 39506
rect 14754 39454 14756 39506
rect 14700 38724 14756 39454
rect 15372 39060 15428 39070
rect 15484 39060 15540 39566
rect 15372 39058 15540 39060
rect 15372 39006 15374 39058
rect 15426 39006 15540 39058
rect 15372 39004 15540 39006
rect 15372 38994 15428 39004
rect 14924 38724 14980 38734
rect 14700 38722 14980 38724
rect 14700 38670 14926 38722
rect 14978 38670 14980 38722
rect 14700 38668 14980 38670
rect 12460 37154 12516 37166
rect 12460 37102 12462 37154
rect 12514 37102 12516 37154
rect 12460 35812 12516 37102
rect 12012 35410 12068 35420
rect 12124 35698 12180 35710
rect 12124 35646 12126 35698
rect 12178 35646 12180 35698
rect 12124 35364 12180 35646
rect 12460 35700 12516 35756
rect 13804 37154 13860 37166
rect 13804 37102 13806 37154
rect 13858 37102 13860 37154
rect 12908 35700 12964 35710
rect 12460 35698 12964 35700
rect 12460 35646 12910 35698
rect 12962 35646 12964 35698
rect 12460 35644 12964 35646
rect 12908 35634 12964 35644
rect 13356 35698 13412 35710
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 12124 35298 12180 35308
rect 12236 35586 12292 35598
rect 12236 35534 12238 35586
rect 12290 35534 12292 35586
rect 11900 34402 11956 34412
rect 11340 34302 11342 34354
rect 11394 34302 11396 34354
rect 11340 34290 11396 34302
rect 12236 34244 12292 35534
rect 13356 35588 13412 35646
rect 13580 35588 13636 35598
rect 13356 35522 13412 35532
rect 13468 35586 13636 35588
rect 13468 35534 13582 35586
rect 13634 35534 13636 35586
rect 13468 35532 13636 35534
rect 12796 35476 12852 35486
rect 12460 35364 12516 35374
rect 12460 35026 12516 35308
rect 12460 34974 12462 35026
rect 12514 34974 12516 35026
rect 12460 34962 12516 34974
rect 12236 34178 12292 34188
rect 12012 34132 12068 34142
rect 12012 34038 12068 34076
rect 12572 34130 12628 34142
rect 12572 34078 12574 34130
rect 12626 34078 12628 34130
rect 12572 34020 12628 34078
rect 12684 34132 12740 34142
rect 12684 34038 12740 34076
rect 12572 33954 12628 33964
rect 11228 33572 11284 33582
rect 11228 33122 11284 33516
rect 12796 33236 12852 35420
rect 13020 34132 13076 34142
rect 13468 34132 13524 35532
rect 13580 35522 13636 35532
rect 13580 34244 13636 34254
rect 13580 34150 13636 34188
rect 13020 34130 13524 34132
rect 13020 34078 13022 34130
rect 13074 34078 13524 34130
rect 13020 34076 13524 34078
rect 13020 34066 13076 34076
rect 12908 34020 12964 34030
rect 12908 33458 12964 33964
rect 13804 33572 13860 37102
rect 12908 33406 12910 33458
rect 12962 33406 12964 33458
rect 12908 33394 12964 33406
rect 13692 33516 13860 33572
rect 12796 33180 12964 33236
rect 11228 33070 11230 33122
rect 11282 33070 11284 33122
rect 11228 32116 11284 33070
rect 11788 33124 11844 33134
rect 11228 32060 11620 32116
rect 11340 28756 11396 28766
rect 11340 27074 11396 28700
rect 11452 28642 11508 28654
rect 11452 28590 11454 28642
rect 11506 28590 11508 28642
rect 11452 28532 11508 28590
rect 11452 28466 11508 28476
rect 11564 28308 11620 32060
rect 11788 28866 11844 33068
rect 12684 31892 12740 31902
rect 12684 31890 12852 31892
rect 12684 31838 12686 31890
rect 12738 31838 12852 31890
rect 12684 31836 12852 31838
rect 12684 31826 12740 31836
rect 11788 28814 11790 28866
rect 11842 28814 11844 28866
rect 11788 28802 11844 28814
rect 11900 29538 11956 29550
rect 11900 29486 11902 29538
rect 11954 29486 11956 29538
rect 11900 28868 11956 29486
rect 12124 29426 12180 29438
rect 12124 29374 12126 29426
rect 12178 29374 12180 29426
rect 12124 29092 12180 29374
rect 12684 29316 12740 29326
rect 12684 29222 12740 29260
rect 12124 29026 12180 29036
rect 12796 28980 12852 31836
rect 12908 29652 12964 33180
rect 13692 31892 13748 33516
rect 13692 31798 13748 31836
rect 13804 31778 13860 31790
rect 13804 31726 13806 31778
rect 13858 31726 13860 31778
rect 13132 30884 13188 30894
rect 13804 30884 13860 31726
rect 13132 30882 13860 30884
rect 13132 30830 13134 30882
rect 13186 30830 13860 30882
rect 13132 30828 13860 30830
rect 13132 30818 13188 30828
rect 12908 29558 12964 29596
rect 13020 29316 13076 29326
rect 13020 29222 13076 29260
rect 11900 28812 12292 28868
rect 11900 28756 11956 28812
rect 11900 28690 11956 28700
rect 11340 27022 11342 27074
rect 11394 27022 11396 27074
rect 11340 27010 11396 27022
rect 11452 28252 11620 28308
rect 12012 28642 12068 28654
rect 12012 28590 12014 28642
rect 12066 28590 12068 28642
rect 11228 26850 11284 26862
rect 11228 26798 11230 26850
rect 11282 26798 11284 26850
rect 11228 26292 11284 26798
rect 11228 26226 11284 26236
rect 11340 26290 11396 26302
rect 11340 26238 11342 26290
rect 11394 26238 11396 26290
rect 11340 25396 11396 26238
rect 11340 25330 11396 25340
rect 11004 25228 11172 25284
rect 10444 23604 10500 23614
rect 10220 23492 10276 23502
rect 8988 22542 8990 22594
rect 9042 22542 9044 22594
rect 8316 22372 8372 22382
rect 8316 22278 8372 22316
rect 8764 22370 8820 22382
rect 8764 22318 8766 22370
rect 8818 22318 8820 22370
rect 7980 22260 8036 22270
rect 7980 22166 8036 22204
rect 8764 22260 8820 22318
rect 8988 22372 9044 22542
rect 8988 22306 9044 22316
rect 9212 22652 9604 22708
rect 8764 22194 8820 22204
rect 7420 21588 7476 21644
rect 7420 21522 7476 21532
rect 7196 21410 7252 21420
rect 7756 21140 7812 21150
rect 6636 21026 6804 21028
rect 6636 20974 6638 21026
rect 6690 20974 6804 21026
rect 6636 20972 6804 20974
rect 7644 21084 7756 21140
rect 6636 20962 6692 20972
rect 6524 20916 6580 20926
rect 6412 20914 6580 20916
rect 6412 20862 6526 20914
rect 6578 20862 6580 20914
rect 6412 20860 6580 20862
rect 5964 20690 6020 20702
rect 5964 20638 5966 20690
rect 6018 20638 6020 20690
rect 5740 20580 5796 20590
rect 5964 20580 6020 20638
rect 6412 20580 6468 20860
rect 6524 20850 6580 20860
rect 5740 20486 5796 20524
rect 5852 20524 6468 20580
rect 5852 20242 5908 20524
rect 5852 20190 5854 20242
rect 5906 20190 5908 20242
rect 5852 20178 5908 20190
rect 5628 20020 5684 20030
rect 5628 19926 5684 19964
rect 7084 19796 7140 19806
rect 6972 19740 7084 19796
rect 6076 18564 6132 18574
rect 5516 18562 6132 18564
rect 5516 18510 6078 18562
rect 6130 18510 6132 18562
rect 5516 18508 6132 18510
rect 6076 18498 6132 18508
rect 6860 18564 6916 18574
rect 6636 18452 6692 18462
rect 6636 18338 6692 18396
rect 6636 18286 6638 18338
rect 6690 18286 6692 18338
rect 6636 18274 6692 18286
rect 6748 18450 6804 18462
rect 6748 18398 6750 18450
rect 6802 18398 6804 18450
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5628 17666 5684 17678
rect 5628 17614 5630 17666
rect 5682 17614 5684 17666
rect 2492 17108 2548 17118
rect 2492 16994 2548 17052
rect 2492 16942 2494 16994
rect 2546 16942 2548 16994
rect 2492 16930 2548 16942
rect 1820 16882 1876 16894
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 13746 1876 16830
rect 5068 16884 5124 16894
rect 5068 16882 5236 16884
rect 5068 16830 5070 16882
rect 5122 16830 5236 16882
rect 5068 16828 5236 16830
rect 5068 16818 5124 16828
rect 4620 16772 4676 16782
rect 4620 16770 4900 16772
rect 4620 16718 4622 16770
rect 4674 16718 4900 16770
rect 4620 16716 4900 16718
rect 4620 16706 4676 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16324 4900 16716
rect 4620 16268 4900 16324
rect 4956 16548 5012 16558
rect 4620 16212 4676 16268
rect 4620 16098 4676 16156
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 4620 16034 4676 16046
rect 4956 16098 5012 16492
rect 4956 16046 4958 16098
rect 5010 16046 5012 16098
rect 4956 16034 5012 16046
rect 5180 16100 5236 16828
rect 5628 16548 5684 17614
rect 5628 16482 5684 16492
rect 5852 17666 5908 17678
rect 5852 17614 5854 17666
rect 5906 17614 5908 17666
rect 5852 17444 5908 17614
rect 6188 17668 6244 17678
rect 6188 17574 6244 17612
rect 6524 17554 6580 17566
rect 6524 17502 6526 17554
rect 6578 17502 6580 17554
rect 6524 17444 6580 17502
rect 5852 17388 6580 17444
rect 6636 17442 6692 17454
rect 6636 17390 6638 17442
rect 6690 17390 6692 17442
rect 5404 16212 5460 16222
rect 5292 16100 5348 16110
rect 5180 16044 5292 16100
rect 5068 15988 5124 15998
rect 5068 15894 5124 15932
rect 5180 15764 5236 16044
rect 5292 16034 5348 16044
rect 5068 15708 5236 15764
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4956 13748 5012 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 11394 1876 13694
rect 4620 13692 4956 13748
rect 2492 13636 2548 13646
rect 2268 13634 2548 13636
rect 2268 13582 2494 13634
rect 2546 13582 2548 13634
rect 2268 13580 2548 13582
rect 2268 12850 2324 13580
rect 2492 13570 2548 13580
rect 4620 13634 4676 13692
rect 4956 13654 5012 13692
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 4620 13570 4676 13582
rect 5068 13524 5124 15708
rect 5404 15148 5460 16156
rect 4956 13468 5124 13524
rect 5180 15092 5460 15148
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2604 12964 2660 12974
rect 2604 12870 2660 12908
rect 2268 12798 2270 12850
rect 2322 12798 2324 12850
rect 2268 12786 2324 12798
rect 4844 12740 4900 12750
rect 4956 12740 5012 13468
rect 4844 12738 5012 12740
rect 4844 12686 4846 12738
rect 4898 12686 5012 12738
rect 4844 12684 5012 12686
rect 2492 12068 2548 12078
rect 2492 11506 2548 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 4620 11620 4676 11630
rect 4620 11506 4676 11564
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11442 4676 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 11172 1876 11342
rect 4844 11172 4900 12684
rect 5180 11954 5236 15092
rect 5852 14420 5908 17388
rect 6412 17108 6468 17118
rect 6412 17014 6468 17052
rect 6300 16884 6356 16894
rect 6524 16884 6580 16894
rect 6076 16882 6356 16884
rect 6076 16830 6302 16882
rect 6354 16830 6356 16882
rect 6076 16828 6356 16830
rect 6076 16210 6132 16828
rect 6300 16818 6356 16828
rect 6412 16882 6580 16884
rect 6412 16830 6526 16882
rect 6578 16830 6580 16882
rect 6412 16828 6580 16830
rect 6300 16548 6356 16558
rect 6076 16158 6078 16210
rect 6130 16158 6132 16210
rect 6076 16146 6132 16158
rect 6188 16212 6244 16222
rect 6188 16098 6244 16156
rect 6188 16046 6190 16098
rect 6242 16046 6244 16098
rect 6188 16034 6244 16046
rect 5964 15988 6020 15998
rect 5964 15426 6020 15932
rect 6300 15764 6356 16492
rect 6188 15708 6356 15764
rect 5964 15374 5966 15426
rect 6018 15374 6020 15426
rect 5964 15362 6020 15374
rect 6076 15428 6132 15438
rect 6076 15334 6132 15372
rect 6188 15148 6244 15708
rect 6300 15540 6356 15550
rect 6412 15540 6468 16828
rect 6524 16818 6580 16828
rect 6636 16548 6692 17390
rect 6748 17444 6804 18398
rect 6860 17666 6916 18508
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 6860 17602 6916 17614
rect 6972 17444 7028 19740
rect 7084 19730 7140 19740
rect 7532 19124 7588 19134
rect 7532 18564 7588 19068
rect 7532 18450 7588 18508
rect 7532 18398 7534 18450
rect 7586 18398 7588 18450
rect 7532 18386 7588 18398
rect 7196 18228 7252 18238
rect 7084 17444 7140 17454
rect 6972 17442 7140 17444
rect 6972 17390 7086 17442
rect 7138 17390 7140 17442
rect 6972 17388 7140 17390
rect 6748 17220 6804 17388
rect 6748 17164 7028 17220
rect 6860 16884 6916 16894
rect 6860 16658 6916 16828
rect 6860 16606 6862 16658
rect 6914 16606 6916 16658
rect 6860 16594 6916 16606
rect 6636 16482 6692 16492
rect 6972 16436 7028 17164
rect 7084 16882 7140 17388
rect 7084 16830 7086 16882
rect 7138 16830 7140 16882
rect 7084 16818 7140 16830
rect 6748 16380 7028 16436
rect 6748 16324 6804 16380
rect 6636 16268 6804 16324
rect 6300 15538 6468 15540
rect 6300 15486 6302 15538
rect 6354 15486 6468 15538
rect 6300 15484 6468 15486
rect 6524 15986 6580 15998
rect 6524 15934 6526 15986
rect 6578 15934 6580 15986
rect 6524 15540 6580 15934
rect 6300 15474 6356 15484
rect 6524 15474 6580 15484
rect 6636 15986 6692 16268
rect 7196 16212 7252 18172
rect 7420 17668 7476 17678
rect 7420 17574 7476 17612
rect 7532 17108 7588 17118
rect 7644 17108 7700 21084
rect 7756 21074 7812 21084
rect 7868 20130 7924 21756
rect 7868 20078 7870 20130
rect 7922 20078 7924 20130
rect 7868 20066 7924 20078
rect 8092 20130 8148 20142
rect 8092 20078 8094 20130
rect 8146 20078 8148 20130
rect 8092 19908 8148 20078
rect 8092 19842 8148 19852
rect 8204 20018 8260 20030
rect 8204 19966 8206 20018
rect 8258 19966 8260 20018
rect 8204 19796 8260 19966
rect 8652 19908 8708 19918
rect 8652 19814 8708 19852
rect 8260 19740 8484 19796
rect 8204 19730 8260 19740
rect 8428 19458 8484 19740
rect 8428 19406 8430 19458
rect 8482 19406 8484 19458
rect 8428 19394 8484 19406
rect 8764 19460 8820 19470
rect 9212 19460 9268 22652
rect 9548 22594 9604 22652
rect 9548 22542 9550 22594
rect 9602 22542 9604 22594
rect 9548 22530 9604 22542
rect 10108 23380 10164 23390
rect 10108 23266 10164 23324
rect 10108 23214 10110 23266
rect 10162 23214 10164 23266
rect 9324 22482 9380 22494
rect 9324 22430 9326 22482
rect 9378 22430 9380 22482
rect 9324 22260 9380 22430
rect 9324 22194 9380 22204
rect 9436 22370 9492 22382
rect 9436 22318 9438 22370
rect 9490 22318 9492 22370
rect 9436 21812 9492 22318
rect 9996 22260 10052 22270
rect 9996 22166 10052 22204
rect 9548 21812 9604 21822
rect 10108 21812 10164 23214
rect 10220 22370 10276 23436
rect 10444 23154 10500 23548
rect 10444 23102 10446 23154
rect 10498 23102 10500 23154
rect 10444 23090 10500 23102
rect 10668 23156 10724 23166
rect 10892 23156 10948 23166
rect 10668 23154 10948 23156
rect 10668 23102 10670 23154
rect 10722 23102 10894 23154
rect 10946 23102 10948 23154
rect 10668 23100 10948 23102
rect 10556 23042 10612 23054
rect 10556 22990 10558 23042
rect 10610 22990 10612 23042
rect 10556 22594 10612 22990
rect 10556 22542 10558 22594
rect 10610 22542 10612 22594
rect 10556 22530 10612 22542
rect 10668 22596 10724 23100
rect 10892 23090 10948 23100
rect 10668 22530 10724 22540
rect 10220 22318 10222 22370
rect 10274 22318 10276 22370
rect 10220 22306 10276 22318
rect 10780 22372 10836 22410
rect 10780 22306 10836 22316
rect 9436 21810 9604 21812
rect 9436 21758 9550 21810
rect 9602 21758 9604 21810
rect 9436 21756 9604 21758
rect 9548 21746 9604 21756
rect 9660 21756 10164 21812
rect 10780 22146 10836 22158
rect 10780 22094 10782 22146
rect 10834 22094 10836 22146
rect 9660 21698 9716 21756
rect 9660 21646 9662 21698
rect 9714 21646 9716 21698
rect 9660 21634 9716 21646
rect 10780 20914 10836 22094
rect 10780 20862 10782 20914
rect 10834 20862 10836 20914
rect 10780 20850 10836 20862
rect 9996 20802 10052 20814
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9660 20580 9716 20590
rect 9996 20580 10052 20750
rect 9660 20578 10052 20580
rect 9660 20526 9662 20578
rect 9714 20526 10052 20578
rect 9660 20524 10052 20526
rect 9660 20244 9716 20524
rect 9884 20356 9940 20366
rect 11004 20356 11060 25228
rect 11340 25172 11396 25182
rect 11340 24724 11396 25116
rect 11452 24946 11508 28252
rect 11676 27076 11732 27086
rect 12012 27076 12068 28590
rect 11676 27074 12068 27076
rect 11676 27022 11678 27074
rect 11730 27022 12068 27074
rect 11676 27020 12068 27022
rect 11676 27010 11732 27020
rect 11900 26852 11956 26862
rect 11564 26850 11956 26852
rect 11564 26798 11902 26850
rect 11954 26798 11956 26850
rect 11564 26796 11956 26798
rect 11564 26290 11620 26796
rect 11900 26786 11956 26796
rect 12012 26850 12068 27020
rect 12236 27074 12292 28812
rect 12236 27022 12238 27074
rect 12290 27022 12292 27074
rect 12236 27010 12292 27022
rect 12460 28532 12516 28542
rect 12460 27074 12516 28476
rect 12796 28530 12852 28924
rect 12908 28868 12964 28878
rect 12908 28642 12964 28812
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12908 28578 12964 28590
rect 12796 28478 12798 28530
rect 12850 28478 12852 28530
rect 12796 28466 12852 28478
rect 12460 27022 12462 27074
rect 12514 27022 12516 27074
rect 12460 27010 12516 27022
rect 12012 26798 12014 26850
rect 12066 26798 12068 26850
rect 12012 26740 12068 26798
rect 12012 26674 12068 26684
rect 12908 26964 12964 26974
rect 11676 26516 11732 26526
rect 11676 26514 12628 26516
rect 11676 26462 11678 26514
rect 11730 26462 12628 26514
rect 11676 26460 12628 26462
rect 11676 26450 11732 26460
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 11564 25956 11620 26238
rect 11788 26290 11844 26302
rect 11788 26238 11790 26290
rect 11842 26238 11844 26290
rect 11788 26180 11844 26238
rect 11788 26114 11844 26124
rect 11900 26290 11956 26302
rect 11900 26238 11902 26290
rect 11954 26238 11956 26290
rect 11564 25890 11620 25900
rect 11900 26068 11956 26238
rect 12348 26292 12404 26302
rect 12348 26198 12404 26236
rect 12572 26290 12628 26460
rect 12908 26402 12964 26908
rect 12908 26350 12910 26402
rect 12962 26350 12964 26402
rect 12908 26338 12964 26350
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12572 26226 12628 26238
rect 11900 25284 11956 26012
rect 12796 26068 12852 26078
rect 13132 26068 13188 26078
rect 12796 26066 13188 26068
rect 12796 26014 12798 26066
rect 12850 26014 13134 26066
rect 13186 26014 13188 26066
rect 12796 26012 13188 26014
rect 12796 26002 12852 26012
rect 13132 26002 13188 26012
rect 11452 24894 11454 24946
rect 11506 24894 11508 24946
rect 11452 24882 11508 24894
rect 11564 25228 11956 25284
rect 12348 25956 12404 25966
rect 11564 24724 11620 25228
rect 11676 24836 11732 24846
rect 11676 24742 11732 24780
rect 12348 24834 12404 25900
rect 13132 24948 13188 24958
rect 13132 24854 13188 24892
rect 12348 24782 12350 24834
rect 12402 24782 12404 24834
rect 12348 24770 12404 24782
rect 11228 24722 11396 24724
rect 11228 24670 11342 24722
rect 11394 24670 11396 24722
rect 11228 24668 11396 24670
rect 11228 23604 11284 24668
rect 11340 24658 11396 24668
rect 11452 24668 11620 24724
rect 11788 24722 11844 24734
rect 11788 24670 11790 24722
rect 11842 24670 11844 24722
rect 11452 23828 11508 24668
rect 11676 24612 11732 24622
rect 11676 24518 11732 24556
rect 11788 23938 11844 24670
rect 12684 24724 12740 24734
rect 12684 24630 12740 24668
rect 13132 24722 13188 24734
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 12796 24612 12852 24622
rect 12796 24518 12852 24556
rect 11788 23886 11790 23938
rect 11842 23886 11844 23938
rect 11564 23828 11620 23838
rect 11452 23826 11620 23828
rect 11452 23774 11566 23826
rect 11618 23774 11620 23826
rect 11452 23772 11620 23774
rect 11228 23378 11284 23548
rect 11228 23326 11230 23378
rect 11282 23326 11284 23378
rect 11228 23314 11284 23326
rect 11340 23492 11396 23502
rect 11340 21140 11396 23436
rect 11452 23380 11508 23390
rect 11452 23286 11508 23324
rect 11564 23268 11620 23772
rect 11564 23202 11620 23212
rect 11564 22932 11620 22942
rect 11564 22838 11620 22876
rect 11788 21812 11844 23886
rect 12908 23380 12964 23390
rect 12684 23268 12740 23278
rect 12684 23174 12740 23212
rect 11340 21074 11396 21084
rect 11676 21756 11844 21812
rect 11900 22372 11956 22382
rect 9660 20178 9716 20188
rect 9772 20300 9884 20356
rect 9548 20130 9604 20142
rect 9548 20078 9550 20130
rect 9602 20078 9604 20130
rect 8764 19458 9268 19460
rect 8764 19406 8766 19458
rect 8818 19406 9268 19458
rect 8764 19404 9268 19406
rect 9324 19908 9380 19918
rect 8764 19394 8820 19404
rect 8652 19010 8708 19022
rect 8652 18958 8654 19010
rect 8706 18958 8708 19010
rect 7980 18562 8036 18574
rect 7980 18510 7982 18562
rect 8034 18510 8036 18562
rect 7980 18452 8036 18510
rect 7980 18386 8036 18396
rect 8316 18452 8372 18462
rect 8316 18358 8372 18396
rect 8652 18340 8708 18958
rect 8540 18338 8708 18340
rect 8540 18286 8654 18338
rect 8706 18286 8708 18338
rect 8540 18284 8708 18286
rect 8316 17444 8372 17454
rect 8316 17350 8372 17388
rect 7532 17106 7700 17108
rect 7532 17054 7534 17106
rect 7586 17054 7700 17106
rect 7532 17052 7700 17054
rect 7532 16884 7588 17052
rect 7532 16818 7588 16828
rect 6636 15934 6638 15986
rect 6690 15934 6692 15986
rect 6188 15092 6356 15148
rect 6188 14530 6244 14542
rect 6188 14478 6190 14530
rect 6242 14478 6244 14530
rect 6188 14420 6244 14478
rect 5404 14364 6244 14420
rect 5292 13858 5348 13870
rect 5292 13806 5294 13858
rect 5346 13806 5348 13858
rect 5292 12516 5348 13806
rect 5292 12450 5348 12460
rect 5404 12066 5460 14364
rect 5852 13972 5908 13982
rect 6300 13972 6356 15092
rect 6412 15092 6468 15102
rect 6412 14754 6468 15036
rect 6412 14702 6414 14754
rect 6466 14702 6468 14754
rect 6412 14690 6468 14702
rect 6636 14756 6692 15934
rect 6860 16156 7252 16212
rect 6860 16098 6916 16156
rect 6860 16046 6862 16098
rect 6914 16046 6916 16098
rect 6860 15092 6916 16046
rect 6860 15026 6916 15036
rect 6636 14662 6692 14700
rect 6748 14418 6804 14430
rect 6748 14366 6750 14418
rect 6802 14366 6804 14418
rect 6748 14196 6804 14366
rect 6748 14140 7140 14196
rect 5852 13970 6356 13972
rect 5852 13918 5854 13970
rect 5906 13918 6356 13970
rect 5852 13916 6356 13918
rect 6636 13972 6692 13982
rect 7084 13972 7140 14140
rect 7308 13972 7364 13982
rect 7084 13970 7364 13972
rect 7084 13918 7310 13970
rect 7362 13918 7364 13970
rect 7084 13916 7364 13918
rect 5852 13906 5908 13916
rect 5628 13748 5684 13786
rect 5628 13682 5684 13692
rect 5964 13522 6020 13534
rect 5964 13470 5966 13522
rect 6018 13470 6020 13522
rect 5740 12516 5796 12526
rect 5516 12180 5572 12190
rect 5516 12178 5684 12180
rect 5516 12126 5518 12178
rect 5570 12126 5684 12178
rect 5516 12124 5684 12126
rect 5516 12114 5572 12124
rect 5404 12014 5406 12066
rect 5458 12014 5460 12066
rect 5404 12002 5460 12014
rect 5180 11902 5182 11954
rect 5234 11902 5236 11954
rect 5180 11508 5236 11902
rect 5404 11508 5460 11518
rect 5180 11452 5404 11508
rect 5404 11442 5460 11452
rect 5628 11282 5684 12124
rect 5740 11394 5796 12460
rect 5964 12290 6020 13470
rect 5964 12238 5966 12290
rect 6018 12238 6020 12290
rect 5964 11844 6020 12238
rect 6412 12178 6468 12190
rect 6412 12126 6414 12178
rect 6466 12126 6468 12178
rect 6076 12068 6132 12078
rect 6412 12068 6468 12126
rect 6636 12178 6692 13916
rect 7308 13906 7364 13916
rect 7420 13972 7476 13982
rect 7420 13878 7476 13916
rect 7532 13860 7588 13870
rect 7532 13766 7588 13804
rect 6636 12126 6638 12178
rect 6690 12126 6692 12178
rect 6636 12114 6692 12126
rect 6860 13412 6916 13422
rect 6860 12404 6916 13356
rect 7644 13412 7700 17052
rect 8428 15316 8484 15326
rect 8540 15316 8596 18284
rect 8652 18274 8708 18284
rect 8764 18562 8820 18574
rect 8764 18510 8766 18562
rect 8818 18510 8820 18562
rect 8764 17780 8820 18510
rect 8988 18452 9044 18462
rect 8988 18358 9044 18396
rect 9100 17780 9156 17790
rect 8652 17724 9100 17780
rect 8652 17666 8708 17724
rect 9100 17686 9156 17724
rect 8652 17614 8654 17666
rect 8706 17614 8708 17666
rect 8652 17602 8708 17614
rect 8428 15314 8596 15316
rect 8428 15262 8430 15314
rect 8482 15262 8596 15314
rect 8428 15260 8596 15262
rect 8428 15250 8484 15260
rect 8092 15092 8148 15102
rect 8092 14530 8148 15036
rect 8092 14478 8094 14530
rect 8146 14478 8148 14530
rect 8092 14466 8148 14478
rect 8316 14756 8372 14766
rect 8316 14530 8372 14700
rect 8316 14478 8318 14530
rect 8370 14478 8372 14530
rect 8316 14466 8372 14478
rect 8204 14308 8260 14318
rect 8204 14214 8260 14252
rect 7980 13748 8036 13758
rect 8092 13748 8148 13758
rect 7980 13746 8092 13748
rect 7980 13694 7982 13746
rect 8034 13694 8092 13746
rect 7980 13692 8092 13694
rect 7980 13682 8036 13692
rect 7644 13346 7700 13356
rect 8092 12740 8148 13692
rect 8204 13522 8260 13534
rect 8204 13470 8206 13522
rect 8258 13470 8260 13522
rect 8204 12964 8260 13470
rect 8204 12898 8260 12908
rect 8540 12962 8596 15260
rect 8652 15428 8708 15438
rect 8652 15148 8708 15372
rect 9324 15148 9380 19852
rect 9548 19348 9604 20078
rect 9548 15148 9604 19292
rect 9772 18452 9828 20300
rect 9884 20290 9940 20300
rect 10780 20300 11060 20356
rect 11340 20916 11396 20926
rect 10556 20244 10612 20254
rect 9884 20020 9940 20030
rect 10332 20020 10388 20030
rect 9884 20018 10388 20020
rect 9884 19966 9886 20018
rect 9938 19966 10334 20018
rect 10386 19966 10388 20018
rect 9884 19964 10388 19966
rect 9884 19954 9940 19964
rect 10332 19954 10388 19964
rect 10556 20018 10612 20188
rect 10556 19966 10558 20018
rect 10610 19966 10612 20018
rect 10556 19954 10612 19966
rect 10220 19796 10276 19806
rect 10220 19702 10276 19740
rect 9660 18338 9716 18350
rect 9660 18286 9662 18338
rect 9714 18286 9716 18338
rect 9660 17892 9716 18286
rect 9772 17892 9828 18396
rect 9884 17892 9940 17902
rect 9772 17890 9940 17892
rect 9772 17838 9886 17890
rect 9938 17838 9940 17890
rect 9772 17836 9940 17838
rect 9660 17826 9716 17836
rect 9884 17826 9940 17836
rect 10108 17780 10164 17790
rect 10108 17686 10164 17724
rect 10668 17780 10724 17790
rect 10668 17686 10724 17724
rect 9660 17668 9716 17678
rect 9660 17574 9716 17612
rect 10220 17554 10276 17566
rect 10220 17502 10222 17554
rect 10274 17502 10276 17554
rect 9660 16100 9716 16110
rect 9660 16006 9716 16044
rect 10220 15876 10276 17502
rect 10332 15988 10388 15998
rect 10332 15986 10500 15988
rect 10332 15934 10334 15986
rect 10386 15934 10500 15986
rect 10332 15932 10500 15934
rect 10332 15922 10388 15932
rect 10220 15810 10276 15820
rect 8652 15092 9044 15148
rect 8652 14532 8708 14542
rect 8876 14532 8932 14542
rect 8652 14530 8932 14532
rect 8652 14478 8654 14530
rect 8706 14478 8878 14530
rect 8930 14478 8932 14530
rect 8652 14476 8932 14478
rect 8652 14466 8708 14476
rect 8876 14466 8932 14476
rect 8876 14308 8932 14318
rect 8764 14196 8820 14206
rect 8764 13858 8820 14140
rect 8764 13806 8766 13858
rect 8818 13806 8820 13858
rect 8764 13794 8820 13806
rect 8876 13858 8932 14252
rect 8876 13806 8878 13858
rect 8930 13806 8932 13858
rect 8876 13794 8932 13806
rect 8652 13748 8708 13758
rect 8652 13654 8708 13692
rect 8540 12910 8542 12962
rect 8594 12910 8596 12962
rect 8540 12898 8596 12910
rect 8428 12852 8484 12862
rect 8428 12758 8484 12796
rect 8204 12740 8260 12750
rect 8092 12738 8260 12740
rect 8092 12686 8206 12738
rect 8258 12686 8260 12738
rect 8092 12684 8260 12686
rect 8204 12674 8260 12684
rect 7868 12516 7924 12526
rect 7756 12404 7812 12414
rect 6860 12178 6916 12348
rect 7084 12402 7812 12404
rect 7084 12350 7758 12402
rect 7810 12350 7812 12402
rect 7084 12348 7812 12350
rect 7084 12290 7140 12348
rect 7756 12338 7812 12348
rect 7868 12402 7924 12460
rect 7868 12350 7870 12402
rect 7922 12350 7924 12402
rect 7868 12338 7924 12350
rect 8428 12404 8484 12414
rect 8428 12310 8484 12348
rect 7084 12238 7086 12290
rect 7138 12238 7140 12290
rect 7084 12226 7140 12238
rect 6860 12126 6862 12178
rect 6914 12126 6916 12178
rect 6860 12114 6916 12126
rect 7420 12180 7476 12190
rect 7420 12086 7476 12124
rect 6076 12066 6468 12068
rect 6076 12014 6078 12066
rect 6130 12014 6468 12066
rect 6076 12012 6468 12014
rect 6076 12002 6132 12012
rect 6412 11956 6468 12012
rect 6524 12068 6580 12078
rect 6524 11974 6580 12012
rect 8988 12068 9044 15092
rect 9212 15092 9380 15148
rect 9436 15092 9604 15148
rect 10332 15540 10388 15550
rect 10332 15426 10388 15484
rect 10444 15538 10500 15932
rect 10444 15486 10446 15538
rect 10498 15486 10500 15538
rect 10444 15474 10500 15486
rect 10332 15374 10334 15426
rect 10386 15374 10388 15426
rect 9212 14644 9268 15092
rect 9212 14530 9268 14588
rect 9212 14478 9214 14530
rect 9266 14478 9268 14530
rect 9212 14466 9268 14478
rect 9436 14420 9492 15092
rect 9660 14644 9716 14654
rect 9660 14550 9716 14588
rect 10108 14644 10164 14654
rect 9436 14364 9716 14420
rect 9100 14306 9156 14318
rect 9100 14254 9102 14306
rect 9154 14254 9156 14306
rect 9100 12852 9156 14254
rect 9436 14196 9492 14364
rect 9436 14130 9492 14140
rect 9660 13972 9716 14364
rect 10108 14084 10164 14588
rect 9660 13970 9940 13972
rect 9660 13918 9662 13970
rect 9714 13918 9940 13970
rect 9660 13916 9940 13918
rect 9660 13906 9716 13916
rect 9100 12786 9156 12796
rect 9212 13860 9268 13870
rect 6412 11890 6468 11900
rect 7644 11956 7700 11966
rect 7644 11862 7700 11900
rect 5964 11788 6244 11844
rect 6188 11620 6244 11788
rect 6188 11526 6244 11564
rect 6412 11508 6468 11518
rect 6412 11414 6468 11452
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5740 11330 5796 11342
rect 8876 11394 8932 11406
rect 8876 11342 8878 11394
rect 8930 11342 8932 11394
rect 5628 11230 5630 11282
rect 5682 11230 5684 11282
rect 5068 11172 5124 11182
rect 4844 11116 5068 11172
rect 1820 11106 1876 11116
rect 5068 11078 5124 11116
rect 4284 10500 4340 10510
rect 2156 10388 2212 10398
rect 2156 9938 2212 10332
rect 2156 9886 2158 9938
rect 2210 9886 2212 9938
rect 2156 9874 2212 9886
rect 4284 9938 4340 10444
rect 5628 10498 5684 11230
rect 6300 11284 6356 11294
rect 5740 10612 5796 10622
rect 6076 10612 6132 10622
rect 5740 10610 6132 10612
rect 5740 10558 5742 10610
rect 5794 10558 6078 10610
rect 6130 10558 6132 10610
rect 5740 10556 6132 10558
rect 5740 10546 5796 10556
rect 6076 10546 6132 10556
rect 6300 10610 6356 11228
rect 6524 11172 6580 11182
rect 6524 11170 6692 11172
rect 6524 11118 6526 11170
rect 6578 11118 6692 11170
rect 6524 11116 6692 11118
rect 6524 11106 6580 11116
rect 6300 10558 6302 10610
rect 6354 10558 6356 10610
rect 6300 10546 6356 10558
rect 6636 10610 6692 11116
rect 6636 10558 6638 10610
rect 6690 10558 6692 10610
rect 6636 10546 6692 10558
rect 7084 10612 7140 10622
rect 7084 10518 7140 10556
rect 5628 10446 5630 10498
rect 5682 10446 5684 10498
rect 5628 10388 5684 10446
rect 6188 10500 6244 10510
rect 6188 10406 6244 10444
rect 7420 10498 7476 10510
rect 7420 10446 7422 10498
rect 7474 10446 7476 10498
rect 5628 10322 5684 10332
rect 6524 10388 6580 10398
rect 6524 10294 6580 10332
rect 7420 10388 7476 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4284 9886 4286 9938
rect 4338 9886 4340 9938
rect 4284 9874 4340 9886
rect 5068 9826 5124 9838
rect 5068 9774 5070 9826
rect 5122 9774 5124 9826
rect 5068 9604 5124 9774
rect 5740 9604 5796 9614
rect 5068 9602 5796 9604
rect 5068 9550 5742 9602
rect 5794 9550 5796 9602
rect 5068 9548 5796 9550
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5740 8428 5796 9548
rect 7420 9268 7476 10332
rect 7420 9202 7476 9212
rect 8092 9604 8148 9614
rect 5404 8372 5796 8428
rect 6076 8932 6132 8942
rect 5404 8260 5460 8372
rect 5404 7474 5460 8204
rect 6076 7586 6132 8876
rect 8092 8370 8148 9548
rect 8876 8428 8932 11342
rect 8092 8318 8094 8370
rect 8146 8318 8148 8370
rect 8092 8306 8148 8318
rect 8652 8372 8932 8428
rect 7420 8260 7476 8270
rect 7420 8166 7476 8204
rect 8428 8260 8484 8270
rect 6076 7534 6078 7586
rect 6130 7534 6132 7586
rect 6076 7522 6132 7534
rect 5404 7422 5406 7474
rect 5458 7422 5460 7474
rect 5404 7410 5460 7422
rect 8428 7476 8484 8204
rect 3500 7364 3556 7374
rect 3276 7362 3556 7364
rect 3276 7310 3502 7362
rect 3554 7310 3556 7362
rect 3276 7308 3556 7310
rect 2716 3444 2772 3454
rect 2940 3444 2996 3454
rect 2716 3442 2996 3444
rect 2716 3390 2718 3442
rect 2770 3390 2942 3442
rect 2994 3390 2996 3442
rect 2716 3388 2996 3390
rect 2716 800 2772 3388
rect 2940 3378 2996 3388
rect 3276 3442 3332 7308
rect 3500 7298 3556 7308
rect 8204 7364 8260 7374
rect 8204 7270 8260 7308
rect 3612 7250 3668 7262
rect 3612 7198 3614 7250
rect 3666 7198 3668 7250
rect 3612 6916 3668 7198
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 3612 6850 3668 6860
rect 8428 6692 8484 7420
rect 8540 7364 8596 7374
rect 8540 7270 8596 7308
rect 8652 7252 8708 8372
rect 8876 7252 8932 7262
rect 8652 7250 8932 7252
rect 8652 7198 8654 7250
rect 8706 7198 8878 7250
rect 8930 7198 8932 7250
rect 8652 7196 8932 7198
rect 8652 7186 8708 7196
rect 8876 7186 8932 7196
rect 8876 6692 8932 6702
rect 8988 6692 9044 12012
rect 9100 11620 9156 11630
rect 9212 11620 9268 13804
rect 9100 11618 9268 11620
rect 9100 11566 9102 11618
rect 9154 11566 9268 11618
rect 9100 11564 9268 11566
rect 9324 11620 9380 11630
rect 9100 11554 9156 11564
rect 9324 11526 9380 11564
rect 9772 11172 9828 11182
rect 9548 11170 9828 11172
rect 9548 11118 9774 11170
rect 9826 11118 9828 11170
rect 9548 11116 9828 11118
rect 9548 10722 9604 11116
rect 9772 11106 9828 11116
rect 9884 10948 9940 13916
rect 10108 13970 10164 14028
rect 10108 13918 10110 13970
rect 10162 13918 10164 13970
rect 10108 13906 10164 13918
rect 10332 13860 10388 15374
rect 10556 15428 10612 15438
rect 10556 15334 10612 15372
rect 10780 14308 10836 20300
rect 11340 20244 11396 20860
rect 11116 19908 11172 19918
rect 11340 19908 11396 20188
rect 11116 19906 11396 19908
rect 11116 19854 11118 19906
rect 11170 19854 11396 19906
rect 11116 19852 11396 19854
rect 11116 19842 11172 19852
rect 11676 19346 11732 21756
rect 11900 20580 11956 22316
rect 12908 20914 12964 23324
rect 13020 23156 13076 23194
rect 13020 23090 13076 23100
rect 13020 22930 13076 22942
rect 13020 22878 13022 22930
rect 13074 22878 13076 22930
rect 13020 22484 13076 22878
rect 13020 22418 13076 22428
rect 13132 22372 13188 24670
rect 13244 23044 13300 30828
rect 13692 29652 13748 29662
rect 13468 29426 13524 29438
rect 13468 29374 13470 29426
rect 13522 29374 13524 29426
rect 13356 28868 13412 28878
rect 13356 26908 13412 28812
rect 13468 28756 13524 29374
rect 13468 27076 13524 28700
rect 13692 28754 13748 29596
rect 13692 28702 13694 28754
rect 13746 28702 13748 28754
rect 13692 28690 13748 28702
rect 13916 27748 13972 38668
rect 14252 38612 14420 38668
rect 14140 37154 14196 37166
rect 14140 37102 14142 37154
rect 14194 37102 14196 37154
rect 14140 36820 14196 37102
rect 14140 36754 14196 36764
rect 14028 35588 14084 35598
rect 14028 35494 14084 35532
rect 14140 32004 14196 32014
rect 13916 27682 13972 27692
rect 14028 31948 14140 32004
rect 13468 27074 13972 27076
rect 13468 27022 13470 27074
rect 13522 27022 13972 27074
rect 13468 27020 13972 27022
rect 13468 27010 13524 27020
rect 13356 26852 13524 26908
rect 13356 26178 13412 26190
rect 13356 26126 13358 26178
rect 13410 26126 13412 26178
rect 13356 26066 13412 26126
rect 13356 26014 13358 26066
rect 13410 26014 13412 26066
rect 13356 23492 13412 26014
rect 13468 25060 13524 26852
rect 13468 25004 13636 25060
rect 13580 24836 13636 25004
rect 13580 24742 13636 24780
rect 13468 24724 13524 24734
rect 13468 24630 13524 24668
rect 13916 23940 13972 27020
rect 14028 26908 14084 31948
rect 14140 31938 14196 31948
rect 14140 29316 14196 29326
rect 14140 29222 14196 29260
rect 14252 26964 14308 27002
rect 14028 26852 14196 26908
rect 14252 26898 14308 26908
rect 14364 26908 14420 38612
rect 14924 37266 14980 38668
rect 15820 38668 15876 46510
rect 16156 46674 16212 46686
rect 16156 46622 16158 46674
rect 16210 46622 16212 46674
rect 15932 45668 15988 45678
rect 15932 45574 15988 45612
rect 15932 44322 15988 44334
rect 15932 44270 15934 44322
rect 15986 44270 15988 44322
rect 15932 44212 15988 44270
rect 15932 44146 15988 44156
rect 16044 44210 16100 44222
rect 16044 44158 16046 44210
rect 16098 44158 16100 44210
rect 16044 43652 16100 44158
rect 16156 44100 16212 46622
rect 16380 46676 16436 46686
rect 16380 46582 16436 46620
rect 16604 46674 16660 46686
rect 16604 46622 16606 46674
rect 16658 46622 16660 46674
rect 16268 46564 16324 46574
rect 16268 46470 16324 46508
rect 16604 46228 16660 46622
rect 17500 46676 17556 46686
rect 17500 46582 17556 46620
rect 16268 46172 16660 46228
rect 17388 46450 17444 46462
rect 17388 46398 17390 46450
rect 17442 46398 17444 46450
rect 16268 46114 16324 46172
rect 16268 46062 16270 46114
rect 16322 46062 16324 46114
rect 16268 46050 16324 46062
rect 16380 45892 16436 45902
rect 16828 45892 16884 45902
rect 16380 45890 16884 45892
rect 16380 45838 16382 45890
rect 16434 45838 16830 45890
rect 16882 45838 16884 45890
rect 16380 45836 16884 45838
rect 16380 45826 16436 45836
rect 16828 45826 16884 45836
rect 16940 45892 16996 45902
rect 16940 45798 16996 45836
rect 17388 45890 17444 46398
rect 17388 45838 17390 45890
rect 17442 45838 17444 45890
rect 17388 45826 17444 45838
rect 17948 45892 18004 45902
rect 17612 45780 17668 45790
rect 17612 45686 17668 45724
rect 17948 45778 18004 45836
rect 17948 45726 17950 45778
rect 18002 45726 18004 45778
rect 17948 45714 18004 45726
rect 16268 45668 16324 45678
rect 16324 45612 16436 45668
rect 16268 45574 16324 45612
rect 16156 44098 16324 44100
rect 16156 44046 16158 44098
rect 16210 44046 16324 44098
rect 16156 44044 16324 44046
rect 16156 44034 16212 44044
rect 16156 43652 16212 43662
rect 16044 43596 16156 43652
rect 16044 42196 16100 43596
rect 16156 43586 16212 43596
rect 16268 43538 16324 44044
rect 16268 43486 16270 43538
rect 16322 43486 16324 43538
rect 16268 43474 16324 43486
rect 16044 42130 16100 42140
rect 16156 40964 16212 40974
rect 16156 39730 16212 40908
rect 16156 39678 16158 39730
rect 16210 39678 16212 39730
rect 16156 39666 16212 39678
rect 15820 38612 16212 38668
rect 14924 37214 14926 37266
rect 14978 37214 14980 37266
rect 14924 37202 14980 37214
rect 15372 37266 15428 37278
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 15372 36484 15428 37214
rect 16156 37266 16212 38612
rect 16380 37940 16436 45612
rect 16716 45666 16772 45678
rect 16716 45614 16718 45666
rect 16770 45614 16772 45666
rect 16716 45108 16772 45614
rect 17500 45332 17556 45342
rect 17500 45330 17892 45332
rect 17500 45278 17502 45330
rect 17554 45278 17892 45330
rect 17500 45276 17892 45278
rect 17500 45266 17556 45276
rect 17276 45108 17332 45118
rect 16716 45106 17332 45108
rect 16716 45054 17278 45106
rect 17330 45054 17332 45106
rect 16716 45052 17332 45054
rect 16492 44324 16548 44334
rect 16716 44324 16772 45052
rect 17276 45042 17332 45052
rect 17612 45108 17668 45118
rect 17836 45108 17892 45276
rect 17612 45106 17780 45108
rect 17612 45054 17614 45106
rect 17666 45054 17780 45106
rect 17612 45052 17780 45054
rect 17612 45042 17668 45052
rect 16492 44322 16772 44324
rect 16492 44270 16494 44322
rect 16546 44270 16772 44322
rect 16492 44268 16772 44270
rect 17276 44324 17332 44334
rect 16492 44258 16548 44268
rect 17276 44230 17332 44268
rect 17500 44322 17556 44334
rect 17500 44270 17502 44322
rect 17554 44270 17556 44322
rect 16828 44212 16884 44222
rect 16492 44100 16548 44110
rect 16492 43538 16548 44044
rect 16828 44100 16884 44156
rect 17388 44100 17444 44110
rect 16828 44098 16996 44100
rect 16828 44046 16830 44098
rect 16882 44046 16996 44098
rect 16828 44044 16996 44046
rect 16828 44034 16884 44044
rect 16492 43486 16494 43538
rect 16546 43486 16548 43538
rect 16492 43474 16548 43486
rect 16716 43314 16772 43326
rect 16716 43262 16718 43314
rect 16770 43262 16772 43314
rect 16716 43092 16772 43262
rect 16828 43316 16884 43326
rect 16828 43222 16884 43260
rect 16716 43026 16772 43036
rect 16940 42980 16996 44044
rect 17388 44006 17444 44044
rect 17500 43876 17556 44270
rect 17724 44324 17780 45052
rect 17724 44258 17780 44268
rect 17500 43810 17556 43820
rect 17836 44210 17892 45052
rect 17836 44158 17838 44210
rect 17890 44158 17892 44210
rect 17612 43426 17668 43438
rect 17612 43374 17614 43426
rect 17666 43374 17668 43426
rect 17612 43092 17668 43374
rect 17388 43036 17612 43092
rect 17052 42980 17108 42990
rect 16940 42924 17052 42980
rect 17052 42914 17108 42924
rect 17388 38668 17444 43036
rect 17612 43026 17668 43036
rect 17612 42868 17668 42878
rect 17836 42868 17892 44158
rect 17612 42866 17892 42868
rect 17612 42814 17614 42866
rect 17666 42814 17892 42866
rect 17612 42812 17892 42814
rect 17948 43988 18004 43998
rect 16380 37874 16436 37884
rect 17276 38612 17444 38668
rect 17500 39732 17556 39742
rect 16156 37214 16158 37266
rect 16210 37214 16212 37266
rect 16156 37202 16212 37214
rect 16716 37828 16772 37838
rect 15484 37154 15540 37166
rect 16380 37156 16436 37166
rect 15484 37102 15486 37154
rect 15538 37102 15540 37154
rect 15484 36708 15540 37102
rect 15484 36642 15540 36652
rect 16268 37154 16436 37156
rect 16268 37102 16382 37154
rect 16434 37102 16436 37154
rect 16268 37100 16436 37102
rect 15708 36484 15764 36494
rect 15372 36482 15876 36484
rect 15372 36430 15710 36482
rect 15762 36430 15876 36482
rect 15372 36428 15876 36430
rect 15708 36418 15764 36428
rect 15596 35700 15652 35710
rect 15596 35606 15652 35644
rect 15148 35586 15204 35598
rect 15148 35534 15150 35586
rect 15202 35534 15204 35586
rect 15036 34132 15092 34142
rect 15036 34038 15092 34076
rect 14476 33124 14532 33134
rect 14476 31890 14532 33068
rect 14924 32676 14980 32686
rect 14924 32582 14980 32620
rect 15148 32674 15204 35534
rect 15708 34914 15764 34926
rect 15708 34862 15710 34914
rect 15762 34862 15764 34914
rect 15708 34692 15764 34862
rect 15708 34626 15764 34636
rect 15596 34244 15652 34254
rect 15484 34242 15652 34244
rect 15484 34190 15598 34242
rect 15650 34190 15652 34242
rect 15484 34188 15652 34190
rect 15484 33124 15540 34188
rect 15596 34178 15652 34188
rect 15484 33058 15540 33068
rect 15596 34018 15652 34030
rect 15596 33966 15598 34018
rect 15650 33966 15652 34018
rect 15148 32622 15150 32674
rect 15202 32622 15204 32674
rect 15148 32610 15204 32622
rect 15484 32676 15540 32686
rect 15484 32582 15540 32620
rect 14476 31838 14478 31890
rect 14530 31838 14532 31890
rect 14476 31826 14532 31838
rect 15036 32450 15092 32462
rect 15036 32398 15038 32450
rect 15090 32398 15092 32450
rect 15036 31778 15092 32398
rect 15148 32004 15204 32014
rect 15148 31910 15204 31948
rect 15036 31726 15038 31778
rect 15090 31726 15092 31778
rect 15036 31714 15092 31726
rect 15596 31666 15652 33966
rect 15596 31614 15598 31666
rect 15650 31614 15652 31666
rect 15596 31602 15652 31614
rect 15820 30322 15876 36428
rect 16044 35924 16100 35934
rect 16044 35698 16100 35868
rect 16044 35646 16046 35698
rect 16098 35646 16100 35698
rect 16044 35634 16100 35646
rect 16268 33460 16324 37100
rect 16380 37090 16436 37100
rect 16492 36708 16548 36718
rect 16492 36372 16548 36652
rect 16604 36372 16660 36382
rect 16492 36370 16660 36372
rect 16492 36318 16606 36370
rect 16658 36318 16660 36370
rect 16492 36316 16660 36318
rect 16604 36306 16660 36316
rect 16604 35924 16660 35934
rect 16604 35830 16660 35868
rect 16716 35588 16772 37772
rect 16828 37154 16884 37166
rect 16828 37102 16830 37154
rect 16882 37102 16884 37154
rect 16828 36484 16884 37102
rect 17164 36484 17220 36494
rect 16828 36482 17220 36484
rect 16828 36430 17166 36482
rect 17218 36430 17220 36482
rect 16828 36428 17220 36430
rect 17164 36418 17220 36428
rect 16716 35522 16772 35532
rect 16940 35476 16996 35486
rect 15932 32562 15988 32574
rect 15932 32510 15934 32562
rect 15986 32510 15988 32562
rect 15932 31556 15988 32510
rect 16268 32450 16324 33404
rect 16268 32398 16270 32450
rect 16322 32398 16324 32450
rect 16268 32386 16324 32398
rect 16380 33458 16436 33470
rect 16380 33406 16382 33458
rect 16434 33406 16436 33458
rect 15932 31490 15988 31500
rect 16156 31668 16212 31678
rect 15820 30270 15822 30322
rect 15874 30270 15876 30322
rect 15484 30212 15540 30222
rect 15372 30210 15540 30212
rect 15372 30158 15486 30210
rect 15538 30158 15540 30210
rect 15372 30156 15540 30158
rect 14364 26852 14980 26908
rect 13356 23426 13412 23436
rect 13804 23938 13972 23940
rect 13804 23886 13918 23938
rect 13970 23886 13972 23938
rect 13804 23884 13972 23886
rect 13244 22978 13300 22988
rect 13692 22484 13748 22494
rect 13692 22390 13748 22428
rect 13132 22306 13188 22316
rect 13468 22260 13524 22270
rect 13468 22166 13524 22204
rect 12908 20862 12910 20914
rect 12962 20862 12964 20914
rect 12908 20850 12964 20862
rect 13580 21588 13636 21598
rect 13804 21588 13860 23884
rect 13916 23874 13972 23884
rect 14028 22932 14084 22942
rect 13916 22372 13972 22382
rect 13916 22278 13972 22316
rect 14028 22370 14084 22876
rect 14028 22318 14030 22370
rect 14082 22318 14084 22370
rect 14028 22306 14084 22318
rect 14028 22146 14084 22158
rect 14028 22094 14030 22146
rect 14082 22094 14084 22146
rect 14028 21812 14084 22094
rect 14140 22036 14196 26852
rect 14700 24948 14756 24958
rect 14700 24050 14756 24892
rect 14700 23998 14702 24050
rect 14754 23998 14756 24050
rect 14700 23986 14756 23998
rect 14364 23156 14420 23166
rect 14364 22596 14420 23100
rect 14924 23156 14980 26852
rect 15260 26404 15316 26414
rect 15260 26310 15316 26348
rect 14980 23100 15092 23156
rect 14924 23090 14980 23100
rect 14364 22370 14420 22540
rect 14364 22318 14366 22370
rect 14418 22318 14420 22370
rect 14364 22306 14420 22318
rect 14812 22372 14868 22382
rect 14812 22278 14868 22316
rect 14140 21980 14420 22036
rect 14028 21756 14308 21812
rect 14252 21698 14308 21756
rect 14252 21646 14254 21698
rect 14306 21646 14308 21698
rect 14252 21634 14308 21646
rect 13580 21586 13860 21588
rect 13580 21534 13582 21586
rect 13634 21534 13860 21586
rect 13580 21532 13860 21534
rect 11676 19294 11678 19346
rect 11730 19294 11732 19346
rect 11676 19282 11732 19294
rect 11788 20132 11844 20142
rect 11788 19234 11844 20076
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 11788 19170 11844 19182
rect 11452 19124 11508 19134
rect 11452 19030 11508 19068
rect 11116 16884 11172 16894
rect 11116 15314 11172 16828
rect 11900 16884 11956 20524
rect 13020 20132 13076 20142
rect 12572 18452 12628 18462
rect 12572 18358 12628 18396
rect 11900 16818 11956 16828
rect 12908 16324 12964 16334
rect 12460 16212 12516 16222
rect 12796 16212 12852 16222
rect 12460 16210 12852 16212
rect 12460 16158 12462 16210
rect 12514 16158 12798 16210
rect 12850 16158 12852 16210
rect 12460 16156 12852 16158
rect 12460 16146 12516 16156
rect 12796 16146 12852 16156
rect 12908 15874 12964 16268
rect 12908 15822 12910 15874
rect 12962 15822 12964 15874
rect 12908 15428 12964 15822
rect 12908 15362 12964 15372
rect 11116 15262 11118 15314
rect 11170 15262 11172 15314
rect 11116 15250 11172 15262
rect 11228 15316 11284 15326
rect 10556 14252 10836 14308
rect 10892 15090 10948 15102
rect 10892 15038 10894 15090
rect 10946 15038 10948 15090
rect 10444 13860 10500 13870
rect 10332 13858 10500 13860
rect 10332 13806 10446 13858
rect 10498 13806 10500 13858
rect 10332 13804 10500 13806
rect 10332 11284 10388 13804
rect 10444 13794 10500 13804
rect 10332 11218 10388 11228
rect 10556 10948 10612 14252
rect 10780 14084 10836 14094
rect 10780 13074 10836 14028
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 10780 13010 10836 13022
rect 10892 13858 10948 15038
rect 10892 13806 10894 13858
rect 10946 13806 10948 13858
rect 10892 11620 10948 13806
rect 11228 13860 11284 15260
rect 13020 14532 13076 20076
rect 13580 18452 13636 21532
rect 13580 18386 13636 18396
rect 13244 18338 13300 18350
rect 13244 18286 13246 18338
rect 13298 18286 13300 18338
rect 13132 17108 13188 17118
rect 13244 17108 13300 18286
rect 14364 17780 14420 21980
rect 15036 20468 15092 23100
rect 15372 22596 15428 30156
rect 15484 30146 15540 30156
rect 15820 30100 15876 30270
rect 15820 30034 15876 30044
rect 16044 30994 16100 31006
rect 16044 30942 16046 30994
rect 16098 30942 16100 30994
rect 15372 22530 15428 22540
rect 15484 29316 15540 29326
rect 15036 20412 15204 20468
rect 14700 20132 14756 20142
rect 14700 20038 14756 20076
rect 15036 20132 15092 20142
rect 15036 20038 15092 20076
rect 14364 17714 14420 17724
rect 14476 18564 14532 18574
rect 13132 17106 13300 17108
rect 13132 17054 13134 17106
rect 13186 17054 13300 17106
rect 13132 17052 13300 17054
rect 13132 17042 13188 17052
rect 13916 16996 13972 17006
rect 13804 16940 13916 16996
rect 13132 16884 13188 16894
rect 13132 16790 13188 16828
rect 13468 16884 13524 16894
rect 13468 16790 13524 16828
rect 13580 16882 13636 16894
rect 13580 16830 13582 16882
rect 13634 16830 13636 16882
rect 13580 16324 13636 16830
rect 13580 16258 13636 16268
rect 13580 16100 13636 16110
rect 13580 16006 13636 16044
rect 13580 15876 13636 15886
rect 13580 15426 13636 15820
rect 13580 15374 13582 15426
rect 13634 15374 13636 15426
rect 13580 15362 13636 15374
rect 12684 14476 13020 14532
rect 11564 14084 11620 14094
rect 11228 13858 11508 13860
rect 11228 13806 11230 13858
rect 11282 13806 11508 13858
rect 11228 13804 11508 13806
rect 11228 13794 11284 13804
rect 11452 12962 11508 13804
rect 11564 13858 11620 14028
rect 11564 13806 11566 13858
rect 11618 13806 11620 13858
rect 11564 13794 11620 13806
rect 11900 13972 11956 13982
rect 11900 13748 11956 13916
rect 12684 13970 12740 14476
rect 13020 14466 13076 14476
rect 12684 13918 12686 13970
rect 12738 13918 12740 13970
rect 12684 13906 12740 13918
rect 13132 14084 13188 14094
rect 13132 13970 13188 14028
rect 13132 13918 13134 13970
rect 13186 13918 13188 13970
rect 13132 13906 13188 13918
rect 12348 13860 12404 13870
rect 12348 13766 12404 13804
rect 11900 13746 12292 13748
rect 11900 13694 11902 13746
rect 11954 13694 12292 13746
rect 11900 13692 12292 13694
rect 11900 13682 11956 13692
rect 11452 12910 11454 12962
rect 11506 12910 11508 12962
rect 11452 12898 11508 12910
rect 11788 13634 11844 13646
rect 11788 13582 11790 13634
rect 11842 13582 11844 13634
rect 11228 12740 11284 12750
rect 11116 12684 11228 12740
rect 11116 11620 11172 12684
rect 11228 12646 11284 12684
rect 11788 12404 11844 13582
rect 12236 13074 12292 13692
rect 12236 13022 12238 13074
rect 12290 13022 12292 13074
rect 12236 13010 12292 13022
rect 13804 12850 13860 16940
rect 13916 16902 13972 16940
rect 14476 16994 14532 18508
rect 14476 16942 14478 16994
rect 14530 16942 14532 16994
rect 14252 15876 14308 15886
rect 13804 12798 13806 12850
rect 13858 12798 13860 12850
rect 13804 12786 13860 12798
rect 13916 15426 13972 15438
rect 13916 15374 13918 15426
rect 13970 15374 13972 15426
rect 13916 13188 13972 15374
rect 14252 15426 14308 15820
rect 14252 15374 14254 15426
rect 14306 15374 14308 15426
rect 14252 15362 14308 15374
rect 14476 14196 14532 16942
rect 14812 17108 14868 17118
rect 14588 16884 14644 16894
rect 14588 16790 14644 16828
rect 14812 16882 14868 17052
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16818 14868 16830
rect 14924 16660 14980 16670
rect 14588 15428 14644 15438
rect 14924 15428 14980 16604
rect 14588 15426 14980 15428
rect 14588 15374 14590 15426
rect 14642 15374 14980 15426
rect 14588 15372 14980 15374
rect 14588 15316 14644 15372
rect 14588 15250 14644 15260
rect 15148 15148 15204 20412
rect 15372 20130 15428 20142
rect 15372 20078 15374 20130
rect 15426 20078 15428 20130
rect 15372 18564 15428 20078
rect 15484 20020 15540 29260
rect 16044 28420 16100 30942
rect 16156 30210 16212 31612
rect 16380 31220 16436 33406
rect 16716 31778 16772 31790
rect 16716 31726 16718 31778
rect 16770 31726 16772 31778
rect 16604 31668 16660 31678
rect 16604 31574 16660 31612
rect 16436 31164 16660 31220
rect 16380 31154 16436 31164
rect 16492 30996 16548 31006
rect 16380 30884 16436 30894
rect 16380 30790 16436 30828
rect 16492 30882 16548 30940
rect 16492 30830 16494 30882
rect 16546 30830 16548 30882
rect 16492 30818 16548 30830
rect 16156 30158 16158 30210
rect 16210 30158 16212 30210
rect 16156 30146 16212 30158
rect 16268 29314 16324 29326
rect 16268 29262 16270 29314
rect 16322 29262 16324 29314
rect 16268 29092 16324 29262
rect 16268 28644 16324 29036
rect 16492 28756 16548 28766
rect 16604 28756 16660 31164
rect 16716 30996 16772 31726
rect 16716 30930 16772 30940
rect 16940 30884 16996 35420
rect 17276 32788 17332 38612
rect 17500 35028 17556 39676
rect 17612 38668 17668 42812
rect 17948 41300 18004 43932
rect 18060 42866 18116 46844
rect 19292 46806 19348 46844
rect 18732 46676 18788 46686
rect 18508 45780 18564 45790
rect 18508 45686 18564 45724
rect 18732 45106 18788 46620
rect 18732 45054 18734 45106
rect 18786 45054 18788 45106
rect 18732 45042 18788 45054
rect 19292 44324 19348 44334
rect 19292 44230 19348 44268
rect 19404 44100 19460 47180
rect 19628 47234 19796 47236
rect 19628 47182 19742 47234
rect 19794 47182 19796 47234
rect 19628 47180 19796 47182
rect 19628 46788 19684 47180
rect 19740 47170 19796 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 45220 19684 46732
rect 20300 46116 20356 47294
rect 20412 46228 20468 48862
rect 20524 47460 20580 47470
rect 20524 47366 20580 47404
rect 20860 47460 20916 47470
rect 21196 47460 21252 47470
rect 20860 47458 21252 47460
rect 20860 47406 20862 47458
rect 20914 47406 21198 47458
rect 21250 47406 21252 47458
rect 20860 47404 21252 47406
rect 20860 47394 20916 47404
rect 21196 47394 21252 47404
rect 21532 47458 21588 47470
rect 21532 47406 21534 47458
rect 21586 47406 21588 47458
rect 21420 47348 21476 47358
rect 21420 47254 21476 47292
rect 20748 47236 20804 47246
rect 20748 47234 21028 47236
rect 20748 47182 20750 47234
rect 20802 47182 21028 47234
rect 20748 47180 21028 47182
rect 20748 47170 20804 47180
rect 20972 46898 21028 47180
rect 20972 46846 20974 46898
rect 21026 46846 21028 46898
rect 20972 46834 21028 46846
rect 20524 46788 20580 46798
rect 20524 46694 20580 46732
rect 21084 46788 21140 46798
rect 21084 46694 21140 46732
rect 20636 46676 20692 46686
rect 20636 46582 20692 46620
rect 20524 46450 20580 46462
rect 20524 46398 20526 46450
rect 20578 46398 20580 46450
rect 20524 46340 20580 46398
rect 21532 46340 21588 47406
rect 21644 46900 21700 48974
rect 21756 49028 21812 49038
rect 21868 49028 21924 49644
rect 22092 49140 22148 49150
rect 22092 49138 22596 49140
rect 22092 49086 22094 49138
rect 22146 49086 22596 49138
rect 22092 49084 22596 49086
rect 22092 49074 22148 49084
rect 21812 48972 21924 49028
rect 21756 48934 21812 48972
rect 21868 47572 21924 48972
rect 21980 49026 22036 49038
rect 21980 48974 21982 49026
rect 22034 48974 22036 49026
rect 21980 48804 22036 48974
rect 22540 49028 22596 49084
rect 22652 49028 22708 49038
rect 22540 49026 22708 49028
rect 22540 48974 22654 49026
rect 22706 48974 22708 49026
rect 22540 48972 22708 48974
rect 22652 48962 22708 48972
rect 22428 48916 22484 48926
rect 22316 48804 22372 48814
rect 21980 48748 22316 48804
rect 22316 48738 22372 48748
rect 21868 47516 22148 47572
rect 21868 47348 21924 47358
rect 21868 47254 21924 47292
rect 21644 46844 21812 46900
rect 20524 46284 21588 46340
rect 20412 46172 21028 46228
rect 20300 46050 20356 46060
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19964 45220 20020 45230
rect 19628 45218 20020 45220
rect 19628 45166 19966 45218
rect 20018 45166 20020 45218
rect 19628 45164 20020 45166
rect 19516 45108 19572 45118
rect 19516 45014 19572 45052
rect 19852 44884 19908 44894
rect 19852 44790 19908 44828
rect 19740 44772 19796 44782
rect 19740 44322 19796 44716
rect 19740 44270 19742 44322
rect 19794 44270 19796 44322
rect 19740 44258 19796 44270
rect 19964 44322 20020 45164
rect 19964 44270 19966 44322
rect 20018 44270 20020 44322
rect 19964 44258 20020 44270
rect 20076 45220 20132 45230
rect 20076 45106 20132 45164
rect 20076 45054 20078 45106
rect 20130 45054 20132 45106
rect 19292 44044 19460 44100
rect 19852 44210 19908 44222
rect 19852 44158 19854 44210
rect 19906 44158 19908 44210
rect 19852 44100 19908 44158
rect 20076 44100 20132 45054
rect 19852 44044 20132 44100
rect 19068 43764 19124 43774
rect 18060 42814 18062 42866
rect 18114 42814 18116 42866
rect 18060 42532 18116 42814
rect 18956 43316 19012 43326
rect 18844 42532 18900 42542
rect 18116 42476 18228 42532
rect 18060 42466 18116 42476
rect 17724 41188 17780 41198
rect 17948 41188 18004 41244
rect 17724 41186 18004 41188
rect 17724 41134 17726 41186
rect 17778 41134 18004 41186
rect 17724 41132 18004 41134
rect 17724 41122 17780 41132
rect 18060 41076 18116 41086
rect 18060 40982 18116 41020
rect 17836 40962 17892 40974
rect 17836 40910 17838 40962
rect 17890 40910 17892 40962
rect 17836 40404 17892 40910
rect 17836 40338 17892 40348
rect 17836 39732 17892 39742
rect 17836 39058 17892 39676
rect 17836 39006 17838 39058
rect 17890 39006 17892 39058
rect 17836 38994 17892 39006
rect 18172 39732 18228 42476
rect 18284 42530 18900 42532
rect 18284 42478 18846 42530
rect 18898 42478 18900 42530
rect 18284 42476 18900 42478
rect 18284 41186 18340 42476
rect 18844 42466 18900 42476
rect 18956 41412 19012 43260
rect 19068 42642 19124 43708
rect 19180 42756 19236 42766
rect 19180 42662 19236 42700
rect 19068 42590 19070 42642
rect 19122 42590 19124 42642
rect 19068 42578 19124 42590
rect 18844 41356 19012 41412
rect 18284 41134 18286 41186
rect 18338 41134 18340 41186
rect 18284 41122 18340 41134
rect 18732 41188 18788 41198
rect 18732 41094 18788 41132
rect 18508 41076 18564 41086
rect 18508 40982 18564 41020
rect 18620 40964 18676 40974
rect 18620 40870 18676 40908
rect 18172 38834 18228 39676
rect 18396 40404 18452 40414
rect 18396 39730 18452 40348
rect 18396 39678 18398 39730
rect 18450 39678 18452 39730
rect 18396 39666 18452 39678
rect 18172 38782 18174 38834
rect 18226 38782 18228 38834
rect 18172 38770 18228 38782
rect 18844 38668 18900 41356
rect 18956 41186 19012 41198
rect 18956 41134 18958 41186
rect 19010 41134 19012 41186
rect 18956 41076 19012 41134
rect 18956 41010 19012 41020
rect 19180 41074 19236 41086
rect 19180 41022 19182 41074
rect 19234 41022 19236 41074
rect 19180 40626 19236 41022
rect 19180 40574 19182 40626
rect 19234 40574 19236 40626
rect 19180 40562 19236 40574
rect 19068 40404 19124 40414
rect 19068 40310 19124 40348
rect 18956 39732 19012 39742
rect 18956 39638 19012 39676
rect 18956 39396 19012 39406
rect 18956 38946 19012 39340
rect 18956 38894 18958 38946
rect 19010 38894 19012 38946
rect 18956 38882 19012 38894
rect 17612 38612 17892 38668
rect 18844 38612 19236 38668
rect 17836 37266 17892 38612
rect 19180 37490 19236 38612
rect 19180 37438 19182 37490
rect 19234 37438 19236 37490
rect 19180 37426 19236 37438
rect 18172 37380 18228 37390
rect 17836 37214 17838 37266
rect 17890 37214 17892 37266
rect 17836 37202 17892 37214
rect 17948 37268 18004 37278
rect 17836 36932 17892 36942
rect 17836 35698 17892 36876
rect 17948 36594 18004 37212
rect 18172 37156 18228 37324
rect 18956 37378 19012 37390
rect 18956 37326 18958 37378
rect 19010 37326 19012 37378
rect 18844 37268 18900 37278
rect 18844 37174 18900 37212
rect 17948 36542 17950 36594
rect 18002 36542 18004 36594
rect 17948 36530 18004 36542
rect 18060 37154 18228 37156
rect 18060 37102 18174 37154
rect 18226 37102 18228 37154
rect 18060 37100 18228 37102
rect 17836 35646 17838 35698
rect 17890 35646 17892 35698
rect 17836 35634 17892 35646
rect 17500 34934 17556 34972
rect 17388 33346 17444 33358
rect 18060 33348 18116 37100
rect 18172 37090 18228 37100
rect 18284 37156 18340 37166
rect 18508 37156 18564 37166
rect 18172 36820 18228 36830
rect 18172 36370 18228 36764
rect 18284 36482 18340 37100
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36418 18340 36430
rect 18396 37154 18564 37156
rect 18396 37102 18510 37154
rect 18562 37102 18564 37154
rect 18396 37100 18564 37102
rect 18172 36318 18174 36370
rect 18226 36318 18228 36370
rect 18172 36306 18228 36318
rect 18284 35698 18340 35710
rect 18284 35646 18286 35698
rect 18338 35646 18340 35698
rect 17388 33294 17390 33346
rect 17442 33294 17444 33346
rect 17388 33124 17444 33294
rect 17388 33058 17444 33068
rect 17836 33292 18116 33348
rect 18172 34692 18228 34702
rect 17276 32732 17444 32788
rect 16940 30210 16996 30828
rect 16940 30158 16942 30210
rect 16994 30158 16996 30210
rect 16940 30146 16996 30158
rect 17276 30100 17332 30110
rect 17276 29652 17332 30044
rect 17276 29586 17332 29596
rect 16828 29316 16884 29326
rect 16828 29222 16884 29260
rect 16548 28700 16884 28756
rect 16492 28662 16548 28700
rect 16268 28578 16324 28588
rect 16044 28364 16436 28420
rect 16380 27186 16436 28364
rect 16380 27134 16382 27186
rect 16434 27134 16436 27186
rect 16380 26908 16436 27134
rect 15596 26852 16436 26908
rect 16828 27186 16884 28700
rect 16828 27134 16830 27186
rect 16882 27134 16884 27186
rect 16828 26908 16884 27134
rect 17388 26908 17444 32732
rect 17724 31220 17780 31230
rect 17724 31126 17780 31164
rect 17836 30324 17892 33292
rect 17948 33124 18004 33134
rect 18172 33124 18228 34636
rect 18004 33068 18228 33124
rect 17948 33030 18004 33068
rect 18284 30884 18340 35646
rect 18396 35364 18452 37100
rect 18508 37090 18564 37100
rect 18956 36036 19012 37326
rect 18956 35980 19236 36036
rect 18508 35588 18564 35598
rect 18508 35586 18676 35588
rect 18508 35534 18510 35586
rect 18562 35534 18676 35586
rect 18508 35532 18676 35534
rect 18508 35522 18564 35532
rect 18396 35308 18564 35364
rect 18508 34802 18564 35308
rect 18620 34916 18676 35532
rect 19068 34916 19124 34926
rect 18620 34914 19124 34916
rect 18620 34862 19070 34914
rect 19122 34862 19124 34914
rect 18620 34860 19124 34862
rect 19068 34850 19124 34860
rect 18508 34750 18510 34802
rect 18562 34750 18564 34802
rect 18508 34738 18564 34750
rect 19180 34690 19236 35980
rect 19292 35698 19348 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20076 43764 20132 43774
rect 19404 43652 19460 43662
rect 19404 42196 19460 43596
rect 20076 43650 20132 43708
rect 20076 43598 20078 43650
rect 20130 43598 20132 43650
rect 20076 43586 20132 43598
rect 19740 43538 19796 43550
rect 19740 43486 19742 43538
rect 19794 43486 19796 43538
rect 19740 43204 19796 43486
rect 19740 43138 19796 43148
rect 20412 43538 20468 43550
rect 20412 43486 20414 43538
rect 20466 43486 20468 43538
rect 20412 43204 20468 43486
rect 20412 43138 20468 43148
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 42140 19796 42196
rect 19628 41188 19684 41198
rect 19740 41188 19796 42140
rect 20412 41748 20468 41758
rect 19964 41188 20020 41198
rect 19740 41186 20020 41188
rect 19740 41134 19966 41186
rect 20018 41134 20020 41186
rect 19740 41132 20020 41134
rect 19628 40962 19684 41132
rect 19964 41122 20020 41132
rect 20412 41186 20468 41692
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 41122 20468 41134
rect 20524 41298 20580 41310
rect 20524 41246 20526 41298
rect 20578 41246 20580 41298
rect 20524 41188 20580 41246
rect 20524 41122 20580 41132
rect 20636 41300 20692 41310
rect 20636 41186 20692 41244
rect 20636 41134 20638 41186
rect 20690 41134 20692 41186
rect 20636 41122 20692 41134
rect 20188 41076 20244 41086
rect 20188 40982 20244 41020
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19628 40404 19684 40910
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20524 40740 20580 40750
rect 20524 40626 20580 40684
rect 20524 40574 20526 40626
rect 20578 40574 20580 40626
rect 20524 40562 20580 40574
rect 19628 40348 20244 40404
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37380 19684 37390
rect 19628 37286 19684 37324
rect 19852 37156 19908 37166
rect 19852 37062 19908 37100
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19292 35646 19294 35698
rect 19346 35646 19348 35698
rect 19292 35634 19348 35646
rect 19740 35700 19796 35710
rect 19740 35606 19796 35644
rect 19852 35586 19908 35598
rect 19852 35534 19854 35586
rect 19906 35534 19908 35586
rect 19628 34916 19684 34926
rect 19852 34916 19908 35534
rect 19628 34914 19908 34916
rect 19628 34862 19630 34914
rect 19682 34862 19908 34914
rect 19628 34860 19908 34862
rect 19628 34850 19684 34860
rect 20076 34804 20132 34814
rect 19740 34802 20132 34804
rect 19740 34750 20078 34802
rect 20130 34750 20132 34802
rect 19740 34748 20132 34750
rect 19740 34692 19796 34748
rect 20076 34738 20132 34748
rect 19180 34638 19182 34690
rect 19234 34638 19236 34690
rect 19180 34626 19236 34638
rect 19292 34636 19796 34692
rect 18620 34468 18676 34478
rect 18620 34130 18676 34412
rect 19292 34242 19348 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19292 34190 19294 34242
rect 19346 34190 19348 34242
rect 19292 34178 19348 34190
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18620 34066 18676 34078
rect 19180 34130 19236 34142
rect 19180 34078 19182 34130
rect 19234 34078 19236 34130
rect 19180 31668 19236 34078
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32788 20244 40348
rect 20300 40402 20356 40414
rect 20860 40404 20916 40414
rect 20300 40350 20302 40402
rect 20354 40350 20356 40402
rect 20300 40292 20356 40350
rect 20636 40402 20916 40404
rect 20636 40350 20862 40402
rect 20914 40350 20916 40402
rect 20636 40348 20916 40350
rect 20636 40292 20692 40348
rect 20860 40338 20916 40348
rect 20300 40236 20692 40292
rect 20524 38724 20580 40236
rect 20972 39284 21028 46172
rect 21644 46116 21700 46126
rect 21644 46022 21700 46060
rect 21756 45892 21812 46844
rect 21196 45836 21812 45892
rect 21980 45890 22036 45902
rect 21980 45838 21982 45890
rect 22034 45838 22036 45890
rect 21196 43652 21252 45836
rect 21980 45332 22036 45838
rect 21868 45106 21924 45118
rect 21868 45054 21870 45106
rect 21922 45054 21924 45106
rect 21308 44322 21364 44334
rect 21308 44270 21310 44322
rect 21362 44270 21364 44322
rect 21308 43876 21364 44270
rect 21868 44324 21924 45054
rect 21980 44772 22036 45276
rect 22092 45108 22148 47516
rect 22428 47460 22484 48860
rect 22764 48802 22820 48814
rect 22764 48750 22766 48802
rect 22818 48750 22820 48802
rect 22764 47684 22820 48750
rect 22876 48804 22932 50316
rect 22988 49812 23044 49822
rect 22988 49026 23044 49756
rect 23212 49698 23268 50430
rect 23436 50484 23492 50494
rect 23212 49646 23214 49698
rect 23266 49646 23268 49698
rect 23212 49634 23268 49646
rect 23324 49924 23380 49934
rect 23324 49028 23380 49868
rect 22988 48974 22990 49026
rect 23042 48974 23044 49026
rect 22988 48962 23044 48974
rect 23212 48972 23380 49028
rect 23436 49026 23492 50428
rect 23996 50484 24052 50494
rect 23996 50390 24052 50428
rect 24108 50482 24164 50494
rect 24108 50430 24110 50482
rect 24162 50430 24164 50482
rect 23436 48974 23438 49026
rect 23490 48974 23492 49026
rect 22876 48710 22932 48748
rect 22764 47618 22820 47628
rect 22484 47404 22596 47460
rect 22428 47394 22484 47404
rect 22204 45890 22260 45902
rect 22204 45838 22206 45890
rect 22258 45838 22260 45890
rect 22204 45220 22260 45838
rect 22316 45220 22372 45230
rect 22204 45164 22316 45220
rect 22316 45154 22372 45164
rect 22092 45106 22260 45108
rect 22092 45054 22094 45106
rect 22146 45054 22260 45106
rect 22092 45052 22260 45054
rect 22092 45042 22148 45052
rect 21980 44706 22036 44716
rect 22092 44436 22148 44446
rect 22092 44342 22148 44380
rect 21868 44268 22036 44324
rect 21308 43820 21476 43876
rect 21308 43652 21364 43662
rect 21196 43650 21364 43652
rect 21196 43598 21310 43650
rect 21362 43598 21364 43650
rect 21196 43596 21364 43598
rect 21308 42756 21364 43596
rect 21420 43540 21476 43820
rect 21644 43540 21700 43550
rect 21980 43540 22036 44268
rect 22204 44212 22260 45052
rect 22428 44996 22484 45006
rect 22428 44902 22484 44940
rect 22316 44882 22372 44894
rect 22316 44830 22318 44882
rect 22370 44830 22372 44882
rect 22316 44772 22372 44830
rect 22316 44706 22372 44716
rect 22540 44436 22596 47404
rect 23212 46900 23268 48972
rect 23436 48962 23492 48974
rect 23548 50370 23604 50382
rect 23548 50318 23550 50370
rect 23602 50318 23604 50370
rect 23548 49922 23604 50318
rect 23548 49870 23550 49922
rect 23602 49870 23604 49922
rect 23548 49028 23604 49870
rect 23548 48962 23604 48972
rect 23660 49140 23716 49150
rect 23660 49026 23716 49084
rect 23660 48974 23662 49026
rect 23714 48974 23716 49026
rect 23660 48962 23716 48974
rect 23996 49026 24052 49038
rect 23996 48974 23998 49026
rect 24050 48974 24052 49026
rect 23996 48916 24052 48974
rect 23548 48802 23604 48814
rect 23548 48750 23550 48802
rect 23602 48750 23604 48802
rect 23548 48692 23604 48750
rect 23548 48626 23604 48636
rect 22988 46844 23268 46900
rect 23660 48244 23716 48254
rect 22764 46676 22820 46686
rect 22652 45890 22708 45902
rect 22652 45838 22654 45890
rect 22706 45838 22708 45890
rect 22652 45220 22708 45838
rect 22764 45890 22820 46620
rect 22764 45838 22766 45890
rect 22818 45838 22820 45890
rect 22764 45826 22820 45838
rect 22988 45892 23044 46844
rect 23100 46674 23156 46686
rect 23100 46622 23102 46674
rect 23154 46622 23156 46674
rect 23100 46116 23156 46622
rect 23212 46676 23268 46686
rect 23212 46582 23268 46620
rect 23324 46676 23380 46686
rect 23660 46676 23716 48188
rect 23996 46900 24052 48860
rect 24108 48804 24164 50430
rect 24332 50484 24388 50542
rect 26124 50594 26180 50652
rect 26348 50708 26404 50718
rect 26348 50614 26404 50652
rect 29148 50706 29204 50718
rect 29148 50654 29150 50706
rect 29202 50654 29204 50706
rect 26124 50542 26126 50594
rect 26178 50542 26180 50594
rect 26124 50530 26180 50542
rect 26460 50594 26516 50606
rect 26460 50542 26462 50594
rect 26514 50542 26516 50594
rect 24332 50418 24388 50428
rect 26012 50484 26068 50494
rect 26460 50428 26516 50542
rect 25900 49924 25956 49934
rect 25676 49868 25900 49924
rect 25564 49140 25620 49150
rect 25564 49026 25620 49084
rect 25676 49138 25732 49868
rect 25900 49830 25956 49868
rect 26012 49924 26068 50428
rect 26236 50372 26516 50428
rect 26796 50482 26852 50494
rect 26796 50430 26798 50482
rect 26850 50430 26852 50482
rect 26236 50034 26292 50372
rect 26236 49982 26238 50034
rect 26290 49982 26292 50034
rect 26236 49970 26292 49982
rect 26796 50036 26852 50430
rect 29148 50484 29204 50654
rect 31276 50708 31332 50718
rect 31276 50614 31332 50652
rect 29148 50418 29204 50428
rect 32060 50596 32116 50606
rect 32396 50596 32452 51214
rect 41692 51266 41972 51268
rect 41692 51214 41918 51266
rect 41970 51214 41972 51266
rect 41692 51212 41972 51214
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35308 50706 35364 50718
rect 35308 50654 35310 50706
rect 35362 50654 35364 50706
rect 35308 50596 35364 50654
rect 36988 50706 37044 50718
rect 36988 50654 36990 50706
rect 37042 50654 37044 50706
rect 32060 50594 32396 50596
rect 32060 50542 32062 50594
rect 32114 50542 32396 50594
rect 32060 50540 32396 50542
rect 26796 49980 26964 50036
rect 26012 49922 26180 49924
rect 26012 49870 26014 49922
rect 26066 49870 26180 49922
rect 26012 49868 26180 49870
rect 26012 49858 26068 49868
rect 25676 49086 25678 49138
rect 25730 49086 25732 49138
rect 25676 49074 25732 49086
rect 25564 48974 25566 49026
rect 25618 48974 25620 49026
rect 25564 48962 25620 48974
rect 25788 49028 25844 49038
rect 26012 49028 26068 49038
rect 25844 49026 26068 49028
rect 25844 48974 26014 49026
rect 26066 48974 26068 49026
rect 25844 48972 26068 48974
rect 25788 48934 25844 48972
rect 26012 48962 26068 48972
rect 24556 48916 24612 48926
rect 24556 48822 24612 48860
rect 25340 48916 25396 48926
rect 25340 48822 25396 48860
rect 24108 48738 24164 48748
rect 24444 48804 24500 48814
rect 24444 47346 24500 48748
rect 26124 48692 26180 49868
rect 26460 49810 26516 49822
rect 26460 49758 26462 49810
rect 26514 49758 26516 49810
rect 26348 49252 26404 49262
rect 26348 49026 26404 49196
rect 26460 49138 26516 49758
rect 26796 49812 26852 49822
rect 26796 49718 26852 49756
rect 26908 49810 26964 49980
rect 27356 49924 27412 49934
rect 27356 49830 27412 49868
rect 27468 49922 27524 49934
rect 27468 49870 27470 49922
rect 27522 49870 27524 49922
rect 26908 49758 26910 49810
rect 26962 49758 26964 49810
rect 26572 49700 26628 49710
rect 26572 49606 26628 49644
rect 26460 49086 26462 49138
rect 26514 49086 26516 49138
rect 26460 49074 26516 49086
rect 26348 48974 26350 49026
rect 26402 48974 26404 49026
rect 26348 48962 26404 48974
rect 26572 48804 26628 48814
rect 25676 48636 26180 48692
rect 26460 48802 26628 48804
rect 26460 48750 26574 48802
rect 26626 48750 26628 48802
rect 26460 48748 26628 48750
rect 24444 47294 24446 47346
rect 24498 47294 24500 47346
rect 24444 47282 24500 47294
rect 24780 47346 24836 47358
rect 24780 47294 24782 47346
rect 24834 47294 24836 47346
rect 24108 46900 24164 46910
rect 23996 46898 24164 46900
rect 23996 46846 24110 46898
rect 24162 46846 24164 46898
rect 23996 46844 24164 46846
rect 23324 46674 23716 46676
rect 23324 46622 23326 46674
rect 23378 46622 23716 46674
rect 23324 46620 23716 46622
rect 23772 46676 23828 46686
rect 23996 46676 24052 46844
rect 24108 46834 24164 46844
rect 23772 46674 24052 46676
rect 23772 46622 23774 46674
rect 23826 46622 24052 46674
rect 23772 46620 24052 46622
rect 23324 46610 23380 46620
rect 23156 46060 23380 46116
rect 23100 46050 23156 46060
rect 23044 45836 23268 45892
rect 22988 45826 23044 45836
rect 22652 45154 22708 45164
rect 22876 45666 22932 45678
rect 22876 45614 22878 45666
rect 22930 45614 22932 45666
rect 22876 44548 22932 45614
rect 22988 45666 23044 45678
rect 22988 45614 22990 45666
rect 23042 45614 23044 45666
rect 22988 45332 23044 45614
rect 22988 45266 23044 45276
rect 23100 45666 23156 45678
rect 23100 45614 23102 45666
rect 23154 45614 23156 45666
rect 23100 45330 23156 45614
rect 23100 45278 23102 45330
rect 23154 45278 23156 45330
rect 23100 45266 23156 45278
rect 23212 45330 23268 45836
rect 23212 45278 23214 45330
rect 23266 45278 23268 45330
rect 23212 45266 23268 45278
rect 22988 44996 23044 45006
rect 23324 44996 23380 46060
rect 23436 45668 23492 46620
rect 23772 46610 23828 46620
rect 24780 45892 24836 47294
rect 24780 45826 24836 45836
rect 24108 45780 24164 45790
rect 24108 45686 24164 45724
rect 24668 45780 24724 45790
rect 23548 45668 23604 45678
rect 23436 45612 23548 45668
rect 22988 44994 23380 44996
rect 22988 44942 22990 44994
rect 23042 44942 23380 44994
rect 22988 44940 23380 44942
rect 22988 44930 23044 44940
rect 22876 44482 22932 44492
rect 22540 44380 22708 44436
rect 22540 44212 22596 44222
rect 22204 44210 22596 44212
rect 22204 44158 22542 44210
rect 22594 44158 22596 44210
rect 22204 44156 22596 44158
rect 22540 44146 22596 44156
rect 22428 43652 22484 43662
rect 22652 43652 22708 44380
rect 22428 43650 22652 43652
rect 22428 43598 22430 43650
rect 22482 43598 22652 43650
rect 22428 43596 22652 43598
rect 22428 43586 22484 43596
rect 22652 43558 22708 43596
rect 21420 43538 22036 43540
rect 21420 43486 21646 43538
rect 21698 43486 22036 43538
rect 21420 43484 22036 43486
rect 22764 43538 22820 43550
rect 22764 43486 22766 43538
rect 22818 43486 22820 43538
rect 21644 43474 21700 43484
rect 21308 42690 21364 42700
rect 21532 41972 21588 41982
rect 21308 41748 21364 41758
rect 21196 41076 21252 41086
rect 21196 40982 21252 41020
rect 21308 41074 21364 41692
rect 21308 41022 21310 41074
rect 21362 41022 21364 41074
rect 21308 41010 21364 41022
rect 21532 40962 21588 41916
rect 21532 40910 21534 40962
rect 21586 40910 21588 40962
rect 21532 40740 21588 40910
rect 21532 40674 21588 40684
rect 21756 41860 21812 41870
rect 21756 41186 21812 41804
rect 21756 41134 21758 41186
rect 21810 41134 21812 41186
rect 21756 40514 21812 41134
rect 21756 40462 21758 40514
rect 21810 40462 21812 40514
rect 21756 40450 21812 40462
rect 21868 40290 21924 43484
rect 22764 43204 22820 43486
rect 22764 43138 22820 43148
rect 21980 43092 22036 43102
rect 21980 42308 22036 43036
rect 23548 42978 23604 45612
rect 24444 45668 24500 45678
rect 24444 45574 24500 45612
rect 24668 45332 24724 45724
rect 25340 45778 25396 45790
rect 25340 45726 25342 45778
rect 25394 45726 25396 45778
rect 24668 45238 24724 45276
rect 25116 45666 25172 45678
rect 25116 45614 25118 45666
rect 25170 45614 25172 45666
rect 25116 44996 25172 45614
rect 25340 45668 25396 45726
rect 25676 45780 25732 48636
rect 26460 48580 26516 48748
rect 26572 48738 26628 48748
rect 26684 48804 26740 48814
rect 25900 48524 26516 48580
rect 25900 48466 25956 48524
rect 25900 48414 25902 48466
rect 25954 48414 25956 48466
rect 25900 48402 25956 48414
rect 25788 48132 25844 48142
rect 26348 48132 26404 48142
rect 26684 48132 26740 48748
rect 25788 48130 26740 48132
rect 25788 48078 25790 48130
rect 25842 48078 26350 48130
rect 26402 48078 26740 48130
rect 25788 48076 26740 48078
rect 25788 48066 25844 48076
rect 25900 47348 25956 47358
rect 25900 47254 25956 47292
rect 26124 47236 26180 47246
rect 25900 45892 25956 45902
rect 25900 45798 25956 45836
rect 25788 45780 25844 45790
rect 25676 45778 25844 45780
rect 25676 45726 25790 45778
rect 25842 45726 25844 45778
rect 25676 45724 25844 45726
rect 25340 45602 25396 45612
rect 25676 45108 25732 45118
rect 25676 45014 25732 45052
rect 23996 44884 24052 44894
rect 23996 44210 24052 44828
rect 25116 44322 25172 44940
rect 25788 44996 25844 45724
rect 25788 44930 25844 44940
rect 26012 45778 26068 45790
rect 26012 45726 26014 45778
rect 26066 45726 26068 45778
rect 25900 44548 25956 44558
rect 25900 44454 25956 44492
rect 25116 44270 25118 44322
rect 25170 44270 25172 44322
rect 25116 44258 25172 44270
rect 23996 44158 23998 44210
rect 24050 44158 24052 44210
rect 23996 44146 24052 44158
rect 23548 42926 23550 42978
rect 23602 42926 23604 42978
rect 23548 42914 23604 42926
rect 24108 43652 24164 43662
rect 23660 42756 23716 42766
rect 23660 42662 23716 42700
rect 23884 42754 23940 42766
rect 23884 42702 23886 42754
rect 23938 42702 23940 42754
rect 23884 42644 23940 42702
rect 24108 42754 24164 43596
rect 25452 42868 25508 42878
rect 26012 42868 26068 45726
rect 26124 44210 26180 47180
rect 26236 47234 26292 47246
rect 26236 47182 26238 47234
rect 26290 47182 26292 47234
rect 26236 46674 26292 47182
rect 26236 46622 26238 46674
rect 26290 46622 26292 46674
rect 26236 45778 26292 46622
rect 26236 45726 26238 45778
rect 26290 45726 26292 45778
rect 26236 45714 26292 45726
rect 26348 45668 26404 48076
rect 26908 47348 26964 49758
rect 27468 49588 27524 49870
rect 27692 49812 27748 49822
rect 32060 49812 32116 50540
rect 32396 50502 32452 50540
rect 35196 50540 35364 50596
rect 35756 50596 35812 50606
rect 33180 50484 33236 50494
rect 33180 50390 33236 50428
rect 33964 50484 34020 50494
rect 35196 50484 35252 50540
rect 35756 50502 35812 50540
rect 33964 50034 34020 50428
rect 34972 50428 35252 50484
rect 36988 50428 37044 50654
rect 40236 50706 40292 50718
rect 40236 50654 40238 50706
rect 40290 50654 40292 50706
rect 39900 50596 39956 50606
rect 39900 50502 39956 50540
rect 34972 50036 35028 50428
rect 36764 50372 37044 50428
rect 37660 50484 37716 50494
rect 33964 49982 33966 50034
rect 34018 49982 34020 50034
rect 33964 49970 34020 49982
rect 34636 49980 35028 50036
rect 35084 50036 35140 50046
rect 33852 49924 33908 49934
rect 33852 49830 33908 49868
rect 33180 49812 33236 49822
rect 27692 49718 27748 49756
rect 31948 49810 33236 49812
rect 31948 49758 32062 49810
rect 32114 49758 33182 49810
rect 33234 49758 33236 49810
rect 31948 49756 33236 49758
rect 28028 49698 28084 49710
rect 28028 49646 28030 49698
rect 28082 49646 28084 49698
rect 28028 49588 28084 49646
rect 27468 49532 28028 49588
rect 27132 48916 27188 48926
rect 27132 48822 27188 48860
rect 27468 48804 27524 49532
rect 28028 49494 28084 49532
rect 29260 49698 29316 49710
rect 29260 49646 29262 49698
rect 29314 49646 29316 49698
rect 29260 49588 29316 49646
rect 31388 49700 31444 49710
rect 31388 49606 31444 49644
rect 29260 49522 29316 49532
rect 27468 48738 27524 48748
rect 27916 47684 27972 47694
rect 27916 47590 27972 47628
rect 26908 47282 26964 47292
rect 28252 47458 28308 47470
rect 28252 47406 28254 47458
rect 28306 47406 28308 47458
rect 28028 47234 28084 47246
rect 28028 47182 28030 47234
rect 28082 47182 28084 47234
rect 26908 46900 26964 46910
rect 26796 46564 26852 46574
rect 26908 46564 26964 46844
rect 28028 46788 28084 47182
rect 28252 47236 28308 47406
rect 31948 47458 32004 49756
rect 32060 49746 32116 49756
rect 33180 49746 33236 49756
rect 34412 49812 34468 49850
rect 34412 49746 34468 49756
rect 34636 49810 34692 49980
rect 34636 49758 34638 49810
rect 34690 49758 34692 49810
rect 34524 49698 34580 49710
rect 34524 49646 34526 49698
rect 34578 49646 34580 49698
rect 34076 49588 34132 49598
rect 34524 49588 34580 49646
rect 34076 49586 34580 49588
rect 34076 49534 34078 49586
rect 34130 49534 34580 49586
rect 34076 49532 34580 49534
rect 34076 49522 34132 49532
rect 34636 49476 34692 49758
rect 34300 49420 34692 49476
rect 34748 49812 34804 49822
rect 33964 48804 34020 48814
rect 31948 47406 31950 47458
rect 32002 47406 32004 47458
rect 31948 47348 32004 47406
rect 33404 48132 33460 48142
rect 28252 47170 28308 47180
rect 31164 47236 31220 47246
rect 31164 47142 31220 47180
rect 31500 47234 31556 47246
rect 31500 47182 31502 47234
rect 31554 47182 31556 47234
rect 28028 46722 28084 46732
rect 30044 46788 30100 46798
rect 30044 46694 30100 46732
rect 30716 46674 30772 46686
rect 30716 46622 30718 46674
rect 30770 46622 30772 46674
rect 27916 46564 27972 46574
rect 26796 46562 26964 46564
rect 26796 46510 26798 46562
rect 26850 46510 26964 46562
rect 26796 46508 26964 46510
rect 26796 46498 26852 46508
rect 26348 45574 26404 45612
rect 26348 44994 26404 45006
rect 26348 44942 26350 44994
rect 26402 44942 26404 44994
rect 26236 44548 26292 44558
rect 26348 44548 26404 44942
rect 26236 44546 26404 44548
rect 26236 44494 26238 44546
rect 26290 44494 26404 44546
rect 26236 44492 26404 44494
rect 26236 44482 26292 44492
rect 26124 44158 26126 44210
rect 26178 44158 26180 44210
rect 26124 43652 26180 44158
rect 26124 43586 26180 43596
rect 26572 43652 26628 43662
rect 26348 42868 26404 42878
rect 26012 42812 26180 42868
rect 25452 42774 25508 42812
rect 24108 42702 24110 42754
rect 24162 42702 24164 42754
rect 24108 42690 24164 42702
rect 25004 42756 25060 42766
rect 25004 42662 25060 42700
rect 25340 42756 25396 42766
rect 21980 41970 22036 42252
rect 21980 41918 21982 41970
rect 22034 41918 22036 41970
rect 21980 41906 22036 41918
rect 22428 42308 22484 42318
rect 22428 41410 22484 42252
rect 23884 42196 23940 42588
rect 24444 42644 24500 42654
rect 24444 42550 24500 42588
rect 25228 42644 25284 42654
rect 25228 42550 25284 42588
rect 23660 42194 23940 42196
rect 23660 42142 23886 42194
rect 23938 42142 23940 42194
rect 23660 42140 23940 42142
rect 23100 41970 23156 41982
rect 23100 41918 23102 41970
rect 23154 41918 23156 41970
rect 23100 41748 23156 41918
rect 23212 41972 23268 41982
rect 23212 41878 23268 41916
rect 23660 41970 23716 42140
rect 23884 42130 23940 42140
rect 24668 42530 24724 42542
rect 24668 42478 24670 42530
rect 24722 42478 24724 42530
rect 24668 42194 24724 42478
rect 24780 42532 24836 42542
rect 25340 42532 25396 42700
rect 25564 42644 25620 42654
rect 26012 42644 26068 42654
rect 25564 42642 26068 42644
rect 25564 42590 25566 42642
rect 25618 42590 26014 42642
rect 26066 42590 26068 42642
rect 25564 42588 26068 42590
rect 25564 42578 25620 42588
rect 24780 42530 24948 42532
rect 24780 42478 24782 42530
rect 24834 42478 24948 42530
rect 24780 42476 24948 42478
rect 25340 42476 25508 42532
rect 24780 42466 24836 42476
rect 24668 42142 24670 42194
rect 24722 42142 24724 42194
rect 24668 42130 24724 42142
rect 23660 41918 23662 41970
rect 23714 41918 23716 41970
rect 23660 41906 23716 41918
rect 24220 41970 24276 41982
rect 24220 41918 24222 41970
rect 24274 41918 24276 41970
rect 23436 41860 23492 41870
rect 23100 41682 23156 41692
rect 23324 41858 23492 41860
rect 23324 41806 23438 41858
rect 23490 41806 23492 41858
rect 23324 41804 23492 41806
rect 23324 41524 23380 41804
rect 23436 41794 23492 41804
rect 24220 41860 24276 41918
rect 24556 41972 24612 41982
rect 24556 41878 24612 41916
rect 24220 41794 24276 41804
rect 22428 41358 22430 41410
rect 22482 41358 22484 41410
rect 22428 41346 22484 41358
rect 22876 41468 23380 41524
rect 23996 41748 24052 41758
rect 22652 41188 22708 41198
rect 22652 41094 22708 41132
rect 22876 41186 22932 41468
rect 22876 41134 22878 41186
rect 22930 41134 22932 41186
rect 22876 41122 22932 41134
rect 22764 40962 22820 40974
rect 22764 40910 22766 40962
rect 22818 40910 22820 40962
rect 21868 40238 21870 40290
rect 21922 40238 21924 40290
rect 21868 40226 21924 40238
rect 22428 40514 22484 40526
rect 22428 40462 22430 40514
rect 22482 40462 22484 40514
rect 22428 40404 22484 40462
rect 21644 39732 21700 39742
rect 21644 39638 21700 39676
rect 22092 39732 22148 39742
rect 22092 39618 22148 39676
rect 22092 39566 22094 39618
rect 22146 39566 22148 39618
rect 22092 39554 22148 39566
rect 20972 39218 21028 39228
rect 22092 39284 22148 39294
rect 21084 38724 21140 38734
rect 20524 38722 21140 38724
rect 20524 38670 21086 38722
rect 21138 38670 21140 38722
rect 20524 38668 21140 38670
rect 22092 38668 22148 39228
rect 22428 38668 22484 40348
rect 22764 39730 22820 40910
rect 22764 39678 22766 39730
rect 22818 39678 22820 39730
rect 22764 39666 22820 39678
rect 23996 40402 24052 41692
rect 24892 40964 24948 42476
rect 25452 42196 25508 42476
rect 25564 42196 25620 42206
rect 25452 42194 25620 42196
rect 25452 42142 25566 42194
rect 25618 42142 25620 42194
rect 25452 42140 25620 42142
rect 25676 42196 25732 42588
rect 26012 42578 26068 42588
rect 26124 42420 26180 42812
rect 26348 42774 26404 42812
rect 26572 42642 26628 43596
rect 26684 42868 26740 42878
rect 26684 42774 26740 42812
rect 26572 42590 26574 42642
rect 26626 42590 26628 42642
rect 26572 42578 26628 42590
rect 26012 42364 26180 42420
rect 25788 42196 25844 42206
rect 25676 42140 25788 42196
rect 25564 42130 25620 42140
rect 25788 42102 25844 42140
rect 25116 41972 25172 41982
rect 25116 41878 25172 41916
rect 25676 41858 25732 41870
rect 25676 41806 25678 41858
rect 25730 41806 25732 41858
rect 24892 40908 25284 40964
rect 23996 40350 23998 40402
rect 24050 40350 24052 40402
rect 23996 38834 24052 40350
rect 24892 39732 24948 39742
rect 23996 38782 23998 38834
rect 24050 38782 24052 38834
rect 23996 38770 24052 38782
rect 24556 39730 24948 39732
rect 24556 39678 24894 39730
rect 24946 39678 24948 39730
rect 24556 39676 24948 39678
rect 24556 39058 24612 39676
rect 24892 39666 24948 39676
rect 25228 39618 25284 40908
rect 25228 39566 25230 39618
rect 25282 39566 25284 39618
rect 25228 39554 25284 39566
rect 25564 39620 25620 39630
rect 25676 39620 25732 41806
rect 25900 39732 25956 39742
rect 25564 39618 25732 39620
rect 25564 39566 25566 39618
rect 25618 39566 25732 39618
rect 25564 39564 25732 39566
rect 25788 39730 25956 39732
rect 25788 39678 25902 39730
rect 25954 39678 25956 39730
rect 25788 39676 25956 39678
rect 25788 39618 25844 39676
rect 25900 39666 25956 39676
rect 25788 39566 25790 39618
rect 25842 39566 25844 39618
rect 25564 39554 25620 39564
rect 25788 39554 25844 39566
rect 25340 39396 25396 39406
rect 25340 39302 25396 39340
rect 24556 39006 24558 39058
rect 24610 39006 24612 39058
rect 24556 38668 24612 39006
rect 20524 37266 20580 38668
rect 21084 38658 21140 38668
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20524 37202 20580 37214
rect 21980 38612 22148 38668
rect 22316 38612 22484 38668
rect 23548 38612 24612 38668
rect 25452 39060 25508 39070
rect 20748 37156 20804 37166
rect 21420 37156 21476 37166
rect 20748 37154 21476 37156
rect 20748 37102 20750 37154
rect 20802 37102 21422 37154
rect 21474 37102 21476 37154
rect 20748 37100 21476 37102
rect 20748 37090 20804 37100
rect 20412 35700 20468 35710
rect 20412 32900 20468 35644
rect 20524 35028 20580 35038
rect 20524 34356 20580 34972
rect 20524 34354 20916 34356
rect 20524 34302 20526 34354
rect 20578 34302 20916 34354
rect 20524 34300 20916 34302
rect 20524 34290 20580 34300
rect 20860 34130 20916 34300
rect 20860 34078 20862 34130
rect 20914 34078 20916 34130
rect 20860 34066 20916 34078
rect 20412 32844 20692 32900
rect 20188 32732 20580 32788
rect 19180 31602 19236 31612
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20412 31108 20468 31118
rect 20412 31014 20468 31052
rect 17948 30324 18004 30334
rect 17836 30268 17948 30324
rect 17948 30230 18004 30268
rect 18172 30212 18228 30222
rect 18172 30118 18228 30156
rect 17724 29426 17780 29438
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 17724 29316 17780 29374
rect 18284 29426 18340 30828
rect 19404 30324 19460 30334
rect 19404 30210 19460 30268
rect 19404 30158 19406 30210
rect 19458 30158 19460 30210
rect 19404 30146 19460 30158
rect 18844 30100 18900 30110
rect 18844 30098 19348 30100
rect 18844 30046 18846 30098
rect 18898 30046 19348 30098
rect 18844 30044 19348 30046
rect 18844 30034 18900 30044
rect 18396 29596 18900 29652
rect 18396 29538 18452 29596
rect 18396 29486 18398 29538
rect 18450 29486 18452 29538
rect 18396 29474 18452 29486
rect 18844 29538 18900 29596
rect 18844 29486 18846 29538
rect 18898 29486 18900 29538
rect 18844 29474 18900 29486
rect 18956 29650 19012 29662
rect 18956 29598 18958 29650
rect 19010 29598 19012 29650
rect 18732 29428 18788 29438
rect 18284 29374 18286 29426
rect 18338 29374 18340 29426
rect 18284 29362 18340 29374
rect 18508 29426 18788 29428
rect 18508 29374 18734 29426
rect 18786 29374 18788 29426
rect 18508 29372 18788 29374
rect 17724 29250 17780 29260
rect 17724 29092 17780 29102
rect 17612 28644 17668 28654
rect 17612 28550 17668 28588
rect 16828 26852 17332 26908
rect 17388 26852 17556 26908
rect 15596 26514 15652 26852
rect 15596 26462 15598 26514
rect 15650 26462 15652 26514
rect 15596 26450 15652 26462
rect 16828 24836 16884 24846
rect 16716 24724 16772 24734
rect 15932 22596 15988 22606
rect 15932 22502 15988 22540
rect 16044 22260 16100 22270
rect 16044 22258 16436 22260
rect 16044 22206 16046 22258
rect 16098 22206 16436 22258
rect 16044 22204 16436 22206
rect 16044 22194 16100 22204
rect 16380 21474 16436 22204
rect 16380 21422 16382 21474
rect 16434 21422 16436 21474
rect 16380 21410 16436 21422
rect 16716 20692 16772 24668
rect 16828 24050 16884 24780
rect 17276 24052 17332 26852
rect 16828 23998 16830 24050
rect 16882 23998 16884 24050
rect 16828 23986 16884 23998
rect 16940 24050 17332 24052
rect 16940 23998 17278 24050
rect 17330 23998 17332 24050
rect 16940 23996 17332 23998
rect 16828 21812 16884 21822
rect 16940 21812 16996 23996
rect 17276 23986 17332 23996
rect 16828 21810 16996 21812
rect 16828 21758 16830 21810
rect 16882 21758 16996 21810
rect 16828 21756 16996 21758
rect 16828 21746 16884 21756
rect 16716 20626 16772 20636
rect 16828 21588 16884 21598
rect 16828 20802 16884 21532
rect 17500 21364 17556 26852
rect 17724 26290 17780 29036
rect 18508 28980 18564 29372
rect 18732 29362 18788 29372
rect 18284 28924 18564 28980
rect 18844 29316 18900 29326
rect 18172 28756 18228 28766
rect 18172 28642 18228 28700
rect 18284 28754 18340 28924
rect 18284 28702 18286 28754
rect 18338 28702 18340 28754
rect 18284 28690 18340 28702
rect 18732 28756 18788 28766
rect 18844 28756 18900 29260
rect 18788 28700 18900 28756
rect 18732 28662 18788 28700
rect 18172 28590 18174 28642
rect 18226 28590 18228 28642
rect 18172 28578 18228 28590
rect 18956 26908 19012 29598
rect 19068 27860 19124 27870
rect 19068 27766 19124 27804
rect 18508 26852 19012 26908
rect 17724 26238 17726 26290
rect 17778 26238 17780 26290
rect 17724 26226 17780 26238
rect 18284 26290 18340 26302
rect 18284 26238 18286 26290
rect 18338 26238 18340 26290
rect 18284 26180 18340 26238
rect 18284 26114 18340 26124
rect 18396 26178 18452 26190
rect 18396 26126 18398 26178
rect 18450 26126 18452 26178
rect 18396 25732 18452 26126
rect 18396 25666 18452 25676
rect 17948 25508 18004 25518
rect 17948 25414 18004 25452
rect 18396 25506 18452 25518
rect 18396 25454 18398 25506
rect 18450 25454 18452 25506
rect 18396 25284 18452 25454
rect 18396 25218 18452 25228
rect 18508 24946 18564 26852
rect 18844 26180 18900 26190
rect 18844 26086 18900 26124
rect 19292 25730 19348 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20300 29540 20356 29550
rect 20188 29538 20356 29540
rect 20188 29486 20302 29538
rect 20354 29486 20356 29538
rect 20188 29484 20356 29486
rect 19628 28980 19684 28990
rect 19628 28642 19684 28924
rect 19628 28590 19630 28642
rect 19682 28590 19684 28642
rect 19628 28578 19684 28590
rect 20076 28756 20132 28766
rect 20076 28642 20132 28700
rect 20076 28590 20078 28642
rect 20130 28590 20132 28642
rect 20076 28578 20132 28590
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28084 19684 28094
rect 20188 28084 20244 29484
rect 20300 29474 20356 29484
rect 20412 29426 20468 29438
rect 20412 29374 20414 29426
rect 20466 29374 20468 29426
rect 20300 28756 20356 28766
rect 20412 28756 20468 29374
rect 20300 28754 20468 28756
rect 20300 28702 20302 28754
rect 20354 28702 20468 28754
rect 20300 28700 20468 28702
rect 20300 28690 20356 28700
rect 19628 27858 19684 28028
rect 19740 28028 20244 28084
rect 20300 28084 20356 28094
rect 19740 27970 19796 28028
rect 19740 27918 19742 27970
rect 19794 27918 19796 27970
rect 19740 27906 19796 27918
rect 19628 27806 19630 27858
rect 19682 27806 19684 27858
rect 19628 27794 19684 27806
rect 20188 27860 20244 27870
rect 20300 27860 20356 28028
rect 20188 27858 20356 27860
rect 20188 27806 20190 27858
rect 20242 27806 20356 27858
rect 20188 27804 20356 27806
rect 20188 27794 20244 27804
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19292 25678 19294 25730
rect 19346 25678 19348 25730
rect 19292 25666 19348 25678
rect 19628 25732 19684 25742
rect 19628 25638 19684 25676
rect 18620 25508 18676 25518
rect 18620 25414 18676 25452
rect 19068 25508 19124 25518
rect 19516 25508 19572 25518
rect 19068 25506 19236 25508
rect 19068 25454 19070 25506
rect 19122 25454 19236 25506
rect 19068 25452 19236 25454
rect 19068 25442 19124 25452
rect 18956 25396 19012 25406
rect 18508 24894 18510 24946
rect 18562 24894 18564 24946
rect 18508 24882 18564 24894
rect 18732 25394 19012 25396
rect 18732 25342 18958 25394
rect 19010 25342 19012 25394
rect 18732 25340 19012 25342
rect 18620 24836 18676 24846
rect 18732 24836 18788 25340
rect 18956 25330 19012 25340
rect 19068 25284 19124 25294
rect 18620 24834 18788 24836
rect 18620 24782 18622 24834
rect 18674 24782 18788 24834
rect 18620 24780 18788 24782
rect 18956 24948 19012 24958
rect 18620 24770 18676 24780
rect 18284 24724 18340 24734
rect 18284 24630 18340 24668
rect 18508 23938 18564 23950
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23380 18564 23886
rect 18956 23938 19012 24892
rect 19068 24946 19124 25228
rect 19068 24894 19070 24946
rect 19122 24894 19124 24946
rect 19068 24836 19124 24894
rect 19068 24770 19124 24780
rect 19068 24052 19124 24062
rect 19180 24052 19236 25452
rect 19516 25414 19572 25452
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24948 20244 24958
rect 20076 24612 20132 24622
rect 20188 24612 20244 24892
rect 20076 24610 20244 24612
rect 20076 24558 20078 24610
rect 20130 24558 20244 24610
rect 20076 24556 20244 24558
rect 20076 24546 20132 24556
rect 19068 24050 19236 24052
rect 19068 23998 19070 24050
rect 19122 23998 19236 24050
rect 19068 23996 19236 23998
rect 19068 23986 19124 23996
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23874 19012 23886
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18508 23314 18564 23324
rect 18284 23268 18340 23278
rect 18284 22482 18340 23212
rect 20076 23268 20132 23278
rect 20412 23268 20468 23278
rect 20076 23266 20468 23268
rect 20076 23214 20078 23266
rect 20130 23214 20414 23266
rect 20466 23214 20468 23266
rect 20076 23212 20468 23214
rect 20076 23202 20132 23212
rect 19516 23156 19572 23166
rect 19516 23062 19572 23100
rect 20412 23156 20468 23212
rect 20524 23268 20580 32732
rect 20636 28084 20692 32844
rect 20748 28756 20804 28766
rect 20972 28756 21028 37100
rect 21420 37090 21476 37100
rect 21980 36260 22036 38612
rect 22092 36484 22148 36494
rect 22316 36484 22372 38612
rect 22988 37154 23044 37166
rect 22988 37102 22990 37154
rect 23042 37102 23044 37154
rect 22988 36708 23044 37102
rect 22092 36482 22372 36484
rect 22092 36430 22094 36482
rect 22146 36430 22372 36482
rect 22092 36428 22372 36430
rect 22540 36652 23044 36708
rect 22540 36482 22596 36652
rect 22540 36430 22542 36482
rect 22594 36430 22596 36482
rect 22092 36418 22148 36428
rect 21980 36204 22148 36260
rect 22092 35700 22148 36204
rect 22204 35700 22260 35710
rect 22092 35698 22260 35700
rect 22092 35646 22206 35698
rect 22258 35646 22260 35698
rect 22092 35644 22260 35646
rect 22204 35634 22260 35644
rect 21980 35586 22036 35598
rect 21980 35534 21982 35586
rect 22034 35534 22036 35586
rect 21980 35252 22036 35534
rect 21644 34020 21700 34030
rect 21980 34020 22036 35196
rect 21644 34018 21812 34020
rect 21644 33966 21646 34018
rect 21698 33966 21812 34018
rect 21644 33964 21812 33966
rect 21644 33954 21700 33964
rect 21756 33572 21812 33964
rect 21980 33954 22036 33964
rect 22428 34244 22484 34254
rect 21756 33516 22036 33572
rect 21980 33458 22036 33516
rect 21980 33406 21982 33458
rect 22034 33406 22036 33458
rect 21980 33394 22036 33406
rect 21756 33348 21812 33358
rect 21644 33346 21812 33348
rect 21644 33294 21758 33346
rect 21810 33294 21812 33346
rect 21644 33292 21812 33294
rect 21644 32786 21700 33292
rect 21756 33282 21812 33292
rect 22092 33346 22148 33358
rect 22428 33348 22484 34188
rect 22092 33294 22094 33346
rect 22146 33294 22148 33346
rect 21644 32734 21646 32786
rect 21698 32734 21700 32786
rect 21644 32722 21700 32734
rect 21868 32674 21924 32686
rect 21868 32622 21870 32674
rect 21922 32622 21924 32674
rect 21868 31780 21924 32622
rect 21980 32564 22036 32574
rect 21980 32470 22036 32508
rect 21868 31714 21924 31724
rect 21532 31668 21588 31678
rect 21420 31612 21532 31668
rect 21084 31220 21140 31230
rect 21084 30994 21140 31164
rect 21084 30942 21086 30994
rect 21138 30942 21140 30994
rect 21084 30930 21140 30942
rect 20804 28700 21028 28756
rect 20748 28662 20804 28700
rect 20972 28196 21028 28700
rect 20972 28130 21028 28140
rect 21084 29876 21140 29886
rect 20636 26628 20692 28028
rect 20636 26562 20692 26572
rect 20524 23202 20580 23212
rect 20412 23090 20468 23100
rect 20636 23154 20692 23166
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 18284 22430 18286 22482
rect 18338 22430 18340 22482
rect 18284 22418 18340 22430
rect 18956 22260 19012 22270
rect 18956 22166 19012 22204
rect 20636 22260 20692 23102
rect 17724 22148 17780 22158
rect 17724 21588 17780 22092
rect 18620 22148 18676 22158
rect 18620 22054 18676 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20636 21812 20692 22204
rect 17724 21494 17780 21532
rect 20524 21756 20692 21812
rect 17500 21298 17556 21308
rect 18284 21474 18340 21486
rect 18284 21422 18286 21474
rect 18338 21422 18340 21474
rect 18284 21364 18340 21422
rect 18284 21298 18340 21308
rect 16828 20750 16830 20802
rect 16882 20750 16884 20802
rect 16604 20580 16660 20590
rect 16604 20486 16660 20524
rect 16044 20468 16100 20478
rect 15708 20132 15764 20142
rect 15708 20038 15764 20076
rect 15484 19954 15540 19964
rect 16044 19908 16100 20412
rect 16492 20130 16548 20142
rect 16492 20078 16494 20130
rect 16546 20078 16548 20130
rect 16044 19842 16100 19852
rect 16268 19908 16324 19918
rect 16268 19814 16324 19852
rect 15372 18498 15428 18508
rect 16268 18452 16324 18462
rect 16268 18358 16324 18396
rect 15372 18340 15428 18350
rect 15708 18340 15764 18350
rect 15372 18338 15764 18340
rect 15372 18286 15374 18338
rect 15426 18286 15710 18338
rect 15762 18286 15764 18338
rect 15372 18284 15764 18286
rect 15372 18274 15428 18284
rect 15708 18274 15764 18284
rect 15932 18340 15988 18350
rect 15820 18226 15876 18238
rect 15820 18174 15822 18226
rect 15874 18174 15876 18226
rect 15820 17780 15876 18174
rect 15484 17724 15876 17780
rect 15484 17220 15540 17724
rect 15260 16884 15316 16894
rect 15260 16882 15428 16884
rect 15260 16830 15262 16882
rect 15314 16830 15428 16882
rect 15260 16828 15428 16830
rect 15260 16818 15316 16828
rect 15372 16322 15428 16828
rect 15372 16270 15374 16322
rect 15426 16270 15428 16322
rect 15372 16258 15428 16270
rect 15484 15986 15540 17164
rect 15820 17108 15876 17118
rect 15932 17108 15988 18284
rect 15876 17052 15988 17108
rect 16380 17444 16436 17454
rect 15820 17014 15876 17052
rect 16044 16884 16100 16894
rect 15932 16882 16100 16884
rect 15932 16830 16046 16882
rect 16098 16830 16100 16882
rect 15932 16828 16100 16830
rect 15484 15934 15486 15986
rect 15538 15934 15540 15986
rect 15484 15922 15540 15934
rect 15708 16098 15764 16110
rect 15708 16046 15710 16098
rect 15762 16046 15764 16098
rect 15708 15988 15764 16046
rect 15820 15988 15876 15998
rect 15708 15932 15820 15988
rect 15820 15922 15876 15932
rect 15932 15148 15988 16828
rect 16044 16818 16100 16828
rect 16380 16882 16436 17388
rect 16492 17108 16548 20078
rect 16828 20130 16884 20750
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16828 20066 16884 20078
rect 17500 20018 17556 20030
rect 17500 19966 17502 20018
rect 17554 19966 17556 20018
rect 17500 19908 17556 19966
rect 17052 19348 17108 19358
rect 17052 19254 17108 19292
rect 17052 17444 17108 17454
rect 17052 17350 17108 17388
rect 17500 17444 17556 19852
rect 18172 19906 18228 19918
rect 18172 19854 18174 19906
rect 18226 19854 18228 19906
rect 18172 19348 18228 19854
rect 20300 19906 20356 19918
rect 20300 19854 20302 19906
rect 20354 19854 20356 19906
rect 20300 19684 20356 19854
rect 20300 19618 20356 19628
rect 20524 19796 20580 21756
rect 20636 21586 20692 21598
rect 20636 21534 20638 21586
rect 20690 21534 20692 21586
rect 20636 20020 20692 21534
rect 20748 20020 20804 20030
rect 20636 20018 20916 20020
rect 20636 19966 20750 20018
rect 20802 19966 20916 20018
rect 20636 19964 20916 19966
rect 20748 19954 20804 19964
rect 18172 19282 18228 19292
rect 20412 19460 20468 19470
rect 20188 19012 20244 19022
rect 19628 18956 20188 19012
rect 17836 17666 17892 17678
rect 17836 17614 17838 17666
rect 17890 17614 17892 17666
rect 17836 17444 17892 17614
rect 17500 17442 17892 17444
rect 17500 17390 17502 17442
rect 17554 17390 17892 17442
rect 17500 17388 17892 17390
rect 18620 17554 18676 17566
rect 18620 17502 18622 17554
rect 18674 17502 18676 17554
rect 17500 17220 17556 17388
rect 16492 17042 16548 17052
rect 16716 17164 17556 17220
rect 17612 17220 17668 17230
rect 16380 16830 16382 16882
rect 16434 16830 16436 16882
rect 16380 16818 16436 16830
rect 16604 16882 16660 16894
rect 16604 16830 16606 16882
rect 16658 16830 16660 16882
rect 16156 16772 16212 16782
rect 16156 16678 16212 16716
rect 16492 16660 16548 16670
rect 16492 16566 16548 16604
rect 16604 16324 16660 16830
rect 16604 16258 16660 16268
rect 16716 16100 16772 17164
rect 17388 16994 17444 17006
rect 17388 16942 17390 16994
rect 17442 16942 17444 16994
rect 17276 16884 17332 16894
rect 17388 16884 17444 16942
rect 17612 16994 17668 17164
rect 17612 16942 17614 16994
rect 17666 16942 17668 16994
rect 17612 16930 17668 16942
rect 17948 17108 18004 17118
rect 16716 16034 16772 16044
rect 17164 16828 17276 16884
rect 17332 16828 17444 16884
rect 17500 16884 17556 16894
rect 15148 15092 15316 15148
rect 15148 14532 15204 14542
rect 15148 14438 15204 14476
rect 14476 14140 14980 14196
rect 14364 13860 14420 13870
rect 13468 12740 13524 12750
rect 13524 12684 13748 12740
rect 13468 12646 13524 12684
rect 10892 11564 11060 11620
rect 10668 11284 10724 11294
rect 10668 11190 10724 11228
rect 10892 11282 10948 11294
rect 10892 11230 10894 11282
rect 10946 11230 10948 11282
rect 9548 10670 9550 10722
rect 9602 10670 9604 10722
rect 9548 10658 9604 10670
rect 9772 10892 9940 10948
rect 10444 10892 10612 10948
rect 9660 10498 9716 10510
rect 9660 10446 9662 10498
rect 9714 10446 9716 10498
rect 9660 8932 9716 10446
rect 9660 8866 9716 8876
rect 9772 8428 9828 10892
rect 10332 10836 10388 10846
rect 9996 10834 10388 10836
rect 9996 10782 10334 10834
rect 10386 10782 10388 10834
rect 9996 10780 10388 10782
rect 9884 10724 9940 10734
rect 9996 10724 10052 10780
rect 10332 10770 10388 10780
rect 9884 10722 10052 10724
rect 9884 10670 9886 10722
rect 9938 10670 10052 10722
rect 9884 10668 10052 10670
rect 9884 10658 9940 10668
rect 10108 10612 10164 10622
rect 10444 10612 10500 10892
rect 10892 10836 10948 11230
rect 10108 10610 10500 10612
rect 10108 10558 10110 10610
rect 10162 10558 10500 10610
rect 10108 10556 10500 10558
rect 10108 10546 10164 10556
rect 10444 9938 10500 10556
rect 10444 9886 10446 9938
rect 10498 9886 10500 9938
rect 10444 9874 10500 9886
rect 10556 10780 10948 10836
rect 10556 10722 10612 10780
rect 10556 10670 10558 10722
rect 10610 10670 10612 10722
rect 10556 8428 10612 10670
rect 10668 10612 10724 10622
rect 11004 10612 11060 11564
rect 11116 11526 11172 11564
rect 11452 12348 11844 12404
rect 11452 11394 11508 12348
rect 13580 12178 13636 12190
rect 13580 12126 13582 12178
rect 13634 12126 13636 12178
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 11330 11508 11342
rect 12796 11396 12852 11406
rect 12796 11302 12852 11340
rect 13468 11396 13524 11406
rect 13468 11302 13524 11340
rect 12908 11282 12964 11294
rect 12908 11230 12910 11282
rect 12962 11230 12964 11282
rect 11116 11172 11172 11182
rect 11116 11170 11284 11172
rect 11116 11118 11118 11170
rect 11170 11118 11284 11170
rect 11116 11116 11284 11118
rect 11116 11106 11172 11116
rect 11116 10612 11172 10622
rect 11004 10556 11116 10612
rect 10668 10518 10724 10556
rect 11116 10518 11172 10556
rect 11116 10052 11172 10062
rect 11116 9826 11172 9996
rect 11228 10050 11284 11116
rect 12684 11170 12740 11182
rect 12684 11118 12686 11170
rect 12738 11118 12740 11170
rect 11452 10724 11508 10734
rect 11452 10722 11732 10724
rect 11452 10670 11454 10722
rect 11506 10670 11732 10722
rect 11452 10668 11732 10670
rect 11452 10658 11508 10668
rect 11228 9998 11230 10050
rect 11282 9998 11284 10050
rect 11228 9986 11284 9998
rect 11116 9774 11118 9826
rect 11170 9774 11172 9826
rect 11116 9762 11172 9774
rect 11564 9940 11620 9950
rect 11564 9826 11620 9884
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11564 9762 11620 9774
rect 11676 9828 11732 10668
rect 12460 10500 12516 10510
rect 12348 10052 12404 10062
rect 11788 9828 11844 9838
rect 12348 9828 12404 9996
rect 12460 10050 12516 10444
rect 12460 9998 12462 10050
rect 12514 9998 12516 10050
rect 12460 9986 12516 9998
rect 12684 9940 12740 11118
rect 12908 10724 12964 11230
rect 12908 10658 12964 10668
rect 13468 11170 13524 11182
rect 13468 11118 13470 11170
rect 13522 11118 13524 11170
rect 13468 10500 13524 11118
rect 13468 10434 13524 10444
rect 13580 10498 13636 12126
rect 13692 11618 13748 12684
rect 13916 12178 13972 13132
rect 14140 13412 14196 13422
rect 14140 12290 14196 13356
rect 14140 12238 14142 12290
rect 14194 12238 14196 12290
rect 14140 12226 14196 12238
rect 14364 12290 14420 13804
rect 14588 13412 14644 13422
rect 14588 13074 14644 13356
rect 14588 13022 14590 13074
rect 14642 13022 14644 13074
rect 14588 13010 14644 13022
rect 14364 12238 14366 12290
rect 14418 12238 14420 12290
rect 13916 12126 13918 12178
rect 13970 12126 13972 12178
rect 13916 12114 13972 12126
rect 14252 12066 14308 12078
rect 14252 12014 14254 12066
rect 14306 12014 14308 12066
rect 13692 11566 13694 11618
rect 13746 11566 13748 11618
rect 13692 11554 13748 11566
rect 14028 11620 14084 11630
rect 14028 11394 14084 11564
rect 14252 11508 14308 12014
rect 14028 11342 14030 11394
rect 14082 11342 14084 11394
rect 14028 11330 14084 11342
rect 14140 11452 14308 11508
rect 13580 10446 13582 10498
rect 13634 10446 13636 10498
rect 13580 10434 13636 10446
rect 13692 10722 13748 10734
rect 13692 10670 13694 10722
rect 13746 10670 13748 10722
rect 13692 10052 13748 10670
rect 13916 10724 13972 10734
rect 13916 10630 13972 10668
rect 13580 9996 13748 10052
rect 14028 10052 14084 10062
rect 14140 10052 14196 11452
rect 14252 11284 14308 11294
rect 14364 11284 14420 12238
rect 14252 11282 14420 11284
rect 14252 11230 14254 11282
rect 14306 11230 14420 11282
rect 14252 11228 14420 11230
rect 14924 12290 14980 14140
rect 15148 12740 15204 12750
rect 15148 12402 15204 12684
rect 15260 12628 15316 15092
rect 15372 15092 15988 15148
rect 16044 15988 16100 15998
rect 15372 14420 15428 15092
rect 15708 14532 15764 14542
rect 15708 14438 15764 14476
rect 15372 14326 15428 14364
rect 16044 14308 16100 15932
rect 17164 15764 17220 16828
rect 17276 16818 17332 16828
rect 17388 16324 17444 16334
rect 17388 16210 17444 16268
rect 17388 16158 17390 16210
rect 17442 16158 17444 16210
rect 17388 16146 17444 16158
rect 17276 15988 17332 15998
rect 17276 15894 17332 15932
rect 17500 15988 17556 16828
rect 17948 16882 18004 17052
rect 18172 17108 18228 17118
rect 18620 17108 18676 17502
rect 18172 17106 18676 17108
rect 18172 17054 18174 17106
rect 18226 17054 18676 17106
rect 18172 17052 18676 17054
rect 18172 17042 18228 17052
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17836 16772 17892 16782
rect 17836 16678 17892 16716
rect 17500 15986 17668 15988
rect 17500 15934 17502 15986
rect 17554 15934 17668 15986
rect 17500 15932 17668 15934
rect 17500 15922 17556 15932
rect 17164 15708 17444 15764
rect 17388 15426 17444 15708
rect 17388 15374 17390 15426
rect 17442 15374 17444 15426
rect 17388 15148 17444 15374
rect 17612 15426 17668 15932
rect 17612 15374 17614 15426
rect 17666 15374 17668 15426
rect 17612 15362 17668 15374
rect 17948 15314 18004 16830
rect 19068 16772 19124 16782
rect 18172 15540 18228 15550
rect 18172 15446 18228 15484
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 17388 15092 17556 15148
rect 17388 14532 17444 14542
rect 17388 14438 17444 14476
rect 16044 14214 16100 14252
rect 16380 14420 16436 14430
rect 15932 13188 15988 13198
rect 15932 13094 15988 13132
rect 15596 12964 15652 12974
rect 15260 12562 15316 12572
rect 15484 12962 15652 12964
rect 15484 12910 15598 12962
rect 15650 12910 15652 12962
rect 15484 12908 15652 12910
rect 15148 12350 15150 12402
rect 15202 12350 15204 12402
rect 15148 12338 15204 12350
rect 14924 12238 14926 12290
rect 14978 12238 14980 12290
rect 14252 11218 14308 11228
rect 14924 10724 14980 12238
rect 15148 12068 15204 12078
rect 14924 10658 14980 10668
rect 15036 11620 15092 11630
rect 14028 10050 14196 10052
rect 14028 9998 14030 10050
rect 14082 9998 14196 10050
rect 14028 9996 14196 9998
rect 13244 9940 13300 9950
rect 12740 9884 12852 9940
rect 12684 9874 12740 9884
rect 11676 9772 11788 9828
rect 11788 9734 11844 9772
rect 12236 9826 12404 9828
rect 12236 9774 12350 9826
rect 12402 9774 12404 9826
rect 12236 9772 12404 9774
rect 11004 9604 11060 9614
rect 11004 9510 11060 9548
rect 11228 9604 11284 9614
rect 11228 8428 11284 9548
rect 12124 9604 12180 9614
rect 12124 9510 12180 9548
rect 12124 9268 12180 9278
rect 12236 9268 12292 9772
rect 12348 9762 12404 9772
rect 12684 9716 12740 9726
rect 12684 9622 12740 9660
rect 12124 9266 12292 9268
rect 12124 9214 12126 9266
rect 12178 9214 12292 9266
rect 12124 9212 12292 9214
rect 12124 9202 12180 9212
rect 9772 8372 10052 8428
rect 9100 7250 9156 7262
rect 9100 7198 9102 7250
rect 9154 7198 9156 7250
rect 9100 7140 9156 7198
rect 9100 7084 9268 7140
rect 8428 6690 8820 6692
rect 8428 6638 8430 6690
rect 8482 6638 8820 6690
rect 8428 6636 8820 6638
rect 8428 6626 8484 6636
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 8764 5124 8820 6636
rect 8876 6690 8988 6692
rect 8876 6638 8878 6690
rect 8930 6638 8988 6690
rect 8876 6636 8988 6638
rect 8876 6626 8932 6636
rect 8988 6598 9044 6636
rect 8988 6466 9044 6478
rect 8988 6414 8990 6466
rect 9042 6414 9044 6466
rect 8988 6020 9044 6414
rect 9100 6468 9156 6478
rect 9212 6468 9268 7084
rect 9996 6804 10052 8372
rect 10220 8372 10612 8428
rect 11116 8372 11284 8428
rect 12796 8482 12852 9884
rect 12908 9828 12964 9838
rect 12908 9734 12964 9772
rect 13244 9266 13300 9884
rect 13580 9716 13636 9996
rect 14028 9986 14084 9996
rect 13916 9940 13972 9950
rect 13916 9826 13972 9884
rect 15036 9938 15092 11564
rect 15036 9886 15038 9938
rect 15090 9886 15092 9938
rect 15036 9874 15092 9886
rect 15148 9940 15204 12012
rect 15260 12068 15316 12078
rect 15484 12068 15540 12908
rect 15596 12898 15652 12908
rect 16380 12962 16436 14364
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 16380 12898 16436 12910
rect 17164 14420 17220 14430
rect 17164 12962 17220 14364
rect 17164 12910 17166 12962
rect 17218 12910 17220 12962
rect 17164 12898 17220 12910
rect 17388 13076 17444 13086
rect 17388 12962 17444 13020
rect 17388 12910 17390 12962
rect 17442 12910 17444 12962
rect 17388 12898 17444 12910
rect 16156 12852 16212 12862
rect 16156 12758 16212 12796
rect 16828 12852 16884 12862
rect 16828 12758 16884 12796
rect 15932 12738 15988 12750
rect 15932 12686 15934 12738
rect 15986 12686 15988 12738
rect 15260 12066 15540 12068
rect 15260 12014 15262 12066
rect 15314 12014 15540 12066
rect 15260 12012 15540 12014
rect 15596 12178 15652 12190
rect 15596 12126 15598 12178
rect 15650 12126 15652 12178
rect 15260 12002 15316 12012
rect 15260 11394 15316 11406
rect 15260 11342 15262 11394
rect 15314 11342 15316 11394
rect 15260 10612 15316 11342
rect 15596 10948 15652 12126
rect 15820 12180 15876 12190
rect 15932 12180 15988 12686
rect 16044 12740 16100 12750
rect 16044 12404 16100 12684
rect 16044 12348 16212 12404
rect 16044 12180 16100 12190
rect 15932 12178 16100 12180
rect 15932 12126 16046 12178
rect 16098 12126 16100 12178
rect 15932 12124 16100 12126
rect 15820 12086 15876 12124
rect 16044 12114 16100 12124
rect 15260 10546 15316 10556
rect 15372 10892 15652 10948
rect 15708 12066 15764 12078
rect 15708 12014 15710 12066
rect 15762 12014 15764 12066
rect 13916 9774 13918 9826
rect 13970 9774 13972 9826
rect 13916 9762 13972 9774
rect 14476 9828 14532 9838
rect 14476 9734 14532 9772
rect 13580 9650 13636 9660
rect 14252 9714 14308 9726
rect 14252 9662 14254 9714
rect 14306 9662 14308 9714
rect 13244 9214 13246 9266
rect 13298 9214 13300 9266
rect 13244 9202 13300 9214
rect 14140 9602 14196 9614
rect 14140 9550 14142 9602
rect 14194 9550 14196 9602
rect 12796 8430 12798 8482
rect 12850 8430 12852 8482
rect 12796 8418 12852 8430
rect 14140 8428 14196 9550
rect 14252 9604 14308 9662
rect 14252 9538 14308 9548
rect 14700 9716 14756 9726
rect 14140 8372 14308 8428
rect 10220 8370 10276 8372
rect 10220 8318 10222 8370
rect 10274 8318 10276 8370
rect 10220 8306 10276 8318
rect 10668 8034 10724 8046
rect 10668 7982 10670 8034
rect 10722 7982 10724 8034
rect 10220 7476 10276 7486
rect 10220 7382 10276 7420
rect 10668 7476 10724 7982
rect 11004 7588 11060 7598
rect 11116 7588 11172 8372
rect 12908 8148 12964 8158
rect 12908 8146 13188 8148
rect 12908 8094 12910 8146
rect 12962 8094 13188 8146
rect 12908 8092 13188 8094
rect 12908 8082 12964 8092
rect 11004 7586 11172 7588
rect 11004 7534 11006 7586
rect 11058 7534 11172 7586
rect 11004 7532 11172 7534
rect 11004 7522 11060 7532
rect 10668 6804 10724 7420
rect 13132 7362 13188 8092
rect 13580 7364 13636 7374
rect 13132 7310 13134 7362
rect 13186 7310 13188 7362
rect 13132 7298 13188 7310
rect 13468 7308 13580 7364
rect 9996 6748 10164 6804
rect 9436 6692 9492 6702
rect 9660 6692 9716 6702
rect 9436 6690 9716 6692
rect 9436 6638 9438 6690
rect 9490 6638 9662 6690
rect 9714 6638 9716 6690
rect 9436 6636 9716 6638
rect 9436 6626 9492 6636
rect 9660 6626 9716 6636
rect 9884 6692 9940 6702
rect 9940 6636 10052 6692
rect 9884 6626 9940 6636
rect 9996 6578 10052 6636
rect 9996 6526 9998 6578
rect 10050 6526 10052 6578
rect 9996 6514 10052 6526
rect 9884 6468 9940 6478
rect 9212 6466 9940 6468
rect 9212 6414 9886 6466
rect 9938 6414 9940 6466
rect 9212 6412 9940 6414
rect 9100 6374 9156 6412
rect 9884 6402 9940 6412
rect 10108 6244 10164 6748
rect 10668 6738 10724 6748
rect 12348 6692 12404 6702
rect 10556 6468 10612 6478
rect 9660 6188 10388 6244
rect 9660 6130 9716 6188
rect 9660 6078 9662 6130
rect 9714 6078 9716 6130
rect 9660 6066 9716 6078
rect 10332 6130 10388 6188
rect 10332 6078 10334 6130
rect 10386 6078 10388 6130
rect 10332 6066 10388 6078
rect 9548 6020 9604 6030
rect 8988 6018 9604 6020
rect 8988 5966 9550 6018
rect 9602 5966 9604 6018
rect 8988 5964 9604 5966
rect 9548 5954 9604 5964
rect 9660 5682 9716 5694
rect 9660 5630 9662 5682
rect 9714 5630 9716 5682
rect 9660 5236 9716 5630
rect 9772 5236 9828 5246
rect 9660 5234 9828 5236
rect 9660 5182 9774 5234
rect 9826 5182 9828 5234
rect 9660 5180 9828 5182
rect 9772 5170 9828 5180
rect 10556 5236 10612 6412
rect 10556 5170 10612 5180
rect 11900 5236 11956 5246
rect 11900 5142 11956 5180
rect 12348 5234 12404 6636
rect 13468 6692 13524 7308
rect 13580 7270 13636 7308
rect 13468 6598 13524 6636
rect 14252 6690 14308 8372
rect 14588 8258 14644 8270
rect 14588 8206 14590 8258
rect 14642 8206 14644 8258
rect 14588 7364 14644 8206
rect 14588 7298 14644 7308
rect 14252 6638 14254 6690
rect 14306 6638 14308 6690
rect 14252 6626 14308 6638
rect 14700 6130 14756 9660
rect 15148 9604 15204 9884
rect 15372 9828 15428 10892
rect 15708 10836 15764 12014
rect 15820 11506 15876 11518
rect 15820 11454 15822 11506
rect 15874 11454 15876 11506
rect 15820 11172 15876 11454
rect 15820 11106 15876 11116
rect 15372 9762 15428 9772
rect 15484 10780 15764 10836
rect 15372 9604 15428 9614
rect 15148 9602 15428 9604
rect 15148 9550 15374 9602
rect 15426 9550 15428 9602
rect 15148 9548 15428 9550
rect 15372 9538 15428 9548
rect 15372 8372 15428 8382
rect 15484 8372 15540 10780
rect 15708 10498 15764 10510
rect 15708 10446 15710 10498
rect 15762 10446 15764 10498
rect 15708 9604 15764 10446
rect 16156 9828 16212 12348
rect 16380 12292 16436 12302
rect 16380 12178 16436 12236
rect 17388 12292 17444 12302
rect 17500 12292 17556 15092
rect 17836 15090 17892 15102
rect 17836 15038 17838 15090
rect 17890 15038 17892 15090
rect 17612 14530 17668 14542
rect 17612 14478 17614 14530
rect 17666 14478 17668 14530
rect 17612 13188 17668 14478
rect 17724 14530 17780 14542
rect 17724 14478 17726 14530
rect 17778 14478 17780 14530
rect 17724 14420 17780 14478
rect 17724 14354 17780 14364
rect 17836 14308 17892 15038
rect 17948 14756 18004 15262
rect 18844 15316 18900 15326
rect 18844 15222 18900 15260
rect 17948 14700 18116 14756
rect 17948 14308 18004 14318
rect 17836 14306 18004 14308
rect 17836 14254 17950 14306
rect 18002 14254 18004 14306
rect 17836 14252 18004 14254
rect 17948 14242 18004 14252
rect 17612 13094 17668 13132
rect 17948 13524 18004 13534
rect 17836 12964 17892 12974
rect 17836 12870 17892 12908
rect 17612 12740 17668 12750
rect 17612 12738 17780 12740
rect 17612 12686 17614 12738
rect 17666 12686 17780 12738
rect 17612 12684 17780 12686
rect 17612 12674 17668 12684
rect 17388 12290 17556 12292
rect 17388 12238 17390 12290
rect 17442 12238 17556 12290
rect 17388 12236 17556 12238
rect 17388 12226 17444 12236
rect 16380 12126 16382 12178
rect 16434 12126 16436 12178
rect 16380 12114 16436 12126
rect 17612 12178 17668 12190
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17500 12068 17556 12078
rect 17388 12066 17556 12068
rect 17388 12014 17502 12066
rect 17554 12014 17556 12066
rect 17388 12012 17556 12014
rect 16828 10612 16884 10622
rect 16828 10518 16884 10556
rect 17388 9938 17444 12012
rect 17500 12002 17556 12012
rect 17612 11956 17668 12126
rect 17724 12180 17780 12684
rect 17836 12180 17892 12190
rect 17724 12178 17892 12180
rect 17724 12126 17838 12178
rect 17890 12126 17892 12178
rect 17724 12124 17892 12126
rect 17836 12114 17892 12124
rect 17948 11956 18004 13468
rect 18060 12292 18116 14700
rect 19068 14532 19124 16716
rect 19516 15540 19572 15550
rect 19516 15426 19572 15484
rect 19516 15374 19518 15426
rect 19570 15374 19572 15426
rect 19516 15362 19572 15374
rect 19068 14438 19124 14476
rect 18284 14418 18340 14430
rect 18284 14366 18286 14418
rect 18338 14366 18340 14418
rect 18284 14308 18340 14366
rect 18396 14420 18452 14430
rect 18396 14326 18452 14364
rect 18284 13186 18340 14252
rect 18508 14306 18564 14318
rect 18508 14254 18510 14306
rect 18562 14254 18564 14306
rect 18508 13524 18564 14254
rect 18508 13458 18564 13468
rect 18284 13134 18286 13186
rect 18338 13134 18340 13186
rect 18284 13122 18340 13134
rect 19068 13188 19124 13198
rect 19068 13074 19124 13132
rect 19068 13022 19070 13074
rect 19122 13022 19124 13074
rect 19068 13010 19124 13022
rect 18396 12964 18452 12974
rect 18396 12870 18452 12908
rect 18620 12962 18676 12974
rect 18620 12910 18622 12962
rect 18674 12910 18676 12962
rect 18060 12178 18116 12236
rect 18060 12126 18062 12178
rect 18114 12126 18116 12178
rect 18060 12114 18116 12126
rect 18620 12180 18676 12910
rect 19628 12404 19684 18956
rect 20188 18918 20244 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20300 16996 20356 17006
rect 20188 16994 20356 16996
rect 20188 16942 20302 16994
rect 20354 16942 20356 16994
rect 20188 16940 20356 16942
rect 20076 16884 20132 16894
rect 20076 16790 20132 16828
rect 20188 16882 20244 16940
rect 20300 16930 20356 16940
rect 20188 16830 20190 16882
rect 20242 16830 20244 16882
rect 20188 16818 20244 16830
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20300 15092 20356 15102
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 12404 20020 12414
rect 17612 11900 18004 11956
rect 17724 11732 17780 11742
rect 17724 11508 17780 11676
rect 17500 11506 17780 11508
rect 17500 11454 17726 11506
rect 17778 11454 17780 11506
rect 17500 11452 17780 11454
rect 17500 10834 17556 11452
rect 17724 11442 17780 11452
rect 17500 10782 17502 10834
rect 17554 10782 17556 10834
rect 17500 10612 17556 10782
rect 18620 10836 18676 12124
rect 19516 12402 20020 12404
rect 19516 12350 19966 12402
rect 20018 12350 20020 12402
rect 19516 12348 20020 12350
rect 18732 10836 18788 10846
rect 18620 10834 18788 10836
rect 18620 10782 18734 10834
rect 18786 10782 18788 10834
rect 18620 10780 18788 10782
rect 18732 10770 18788 10780
rect 19516 10612 19572 12348
rect 19964 12338 20020 12348
rect 20300 11620 20356 15036
rect 20300 11554 20356 11564
rect 20412 12066 20468 19404
rect 20524 19234 20580 19740
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19170 20580 19182
rect 20748 17780 20804 17790
rect 20636 17778 20804 17780
rect 20636 17726 20750 17778
rect 20802 17726 20804 17778
rect 20636 17724 20804 17726
rect 20636 16994 20692 17724
rect 20748 17714 20804 17724
rect 20636 16942 20638 16994
rect 20690 16942 20692 16994
rect 20636 16930 20692 16942
rect 20860 16884 20916 19964
rect 20972 16884 21028 16894
rect 20860 16882 21028 16884
rect 20860 16830 20974 16882
rect 21026 16830 21028 16882
rect 20860 16828 21028 16830
rect 20972 15316 21028 16828
rect 21084 16772 21140 29820
rect 21420 29652 21476 31612
rect 21532 31602 21588 31612
rect 22092 31556 22148 33294
rect 21980 31500 22148 31556
rect 22204 33346 22484 33348
rect 22204 33294 22430 33346
rect 22482 33294 22484 33346
rect 22204 33292 22484 33294
rect 21644 31108 21700 31118
rect 21644 31014 21700 31052
rect 21532 30996 21588 31006
rect 21532 30902 21588 30940
rect 21756 30994 21812 31006
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 21756 30212 21812 30942
rect 21980 30434 22036 31500
rect 22092 31108 22148 31118
rect 22204 31108 22260 33292
rect 22428 33282 22484 33292
rect 22540 32788 22596 36430
rect 22876 36484 22932 36494
rect 22652 36372 22708 36382
rect 22652 36278 22708 36316
rect 22876 35810 22932 36428
rect 22876 35758 22878 35810
rect 22930 35758 22932 35810
rect 22876 35746 22932 35758
rect 23100 36482 23156 36494
rect 23100 36430 23102 36482
rect 23154 36430 23156 36482
rect 23100 35476 23156 36430
rect 23548 36482 23604 38612
rect 23996 36596 24052 36606
rect 23996 36594 24612 36596
rect 23996 36542 23998 36594
rect 24050 36542 24612 36594
rect 23996 36540 24612 36542
rect 23996 36530 24052 36540
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 36418 23604 36430
rect 24556 36484 24612 36540
rect 24892 36484 24948 36494
rect 24556 36482 24948 36484
rect 24556 36430 24894 36482
rect 24946 36430 24948 36482
rect 24556 36428 24948 36430
rect 24892 36418 24948 36428
rect 25340 36484 25396 36494
rect 25340 36390 25396 36428
rect 24332 36372 24388 36382
rect 24332 36278 24388 36316
rect 23100 35410 23156 35420
rect 23436 35586 23492 35598
rect 23436 35534 23438 35586
rect 23490 35534 23492 35586
rect 23436 35252 23492 35534
rect 23436 35186 23492 35196
rect 24220 35586 24276 35598
rect 24220 35534 24222 35586
rect 24274 35534 24276 35586
rect 24220 35476 24276 35534
rect 24220 35028 24276 35420
rect 25340 35586 25396 35598
rect 25340 35534 25342 35586
rect 25394 35534 25396 35586
rect 25340 35364 25396 35534
rect 25340 35298 25396 35308
rect 24220 34962 24276 34972
rect 24668 34804 24724 34814
rect 25340 34804 25396 34814
rect 25452 34804 25508 39004
rect 25676 37492 25732 37502
rect 25676 36594 25732 37436
rect 25676 36542 25678 36594
rect 25730 36542 25732 36594
rect 25676 36530 25732 36542
rect 25900 37268 25956 37278
rect 26012 37268 26068 42364
rect 26124 42084 26180 42094
rect 26124 41298 26180 42028
rect 26348 41972 26404 41982
rect 26348 41878 26404 41916
rect 26124 41246 26126 41298
rect 26178 41246 26180 41298
rect 26124 41234 26180 41246
rect 26124 39732 26180 39742
rect 26348 39732 26404 39742
rect 26124 39730 26404 39732
rect 26124 39678 26126 39730
rect 26178 39678 26350 39730
rect 26402 39678 26404 39730
rect 26124 39676 26404 39678
rect 26124 39172 26180 39676
rect 26348 39666 26404 39676
rect 26124 39116 26404 39172
rect 26348 38668 26404 39116
rect 26124 38612 26404 38668
rect 26124 37380 26180 38612
rect 26124 37286 26180 37324
rect 25900 37266 26068 37268
rect 25900 37214 25902 37266
rect 25954 37214 26068 37266
rect 25900 37212 26068 37214
rect 25788 35700 25844 35710
rect 25788 35606 25844 35644
rect 25676 34804 25732 34814
rect 25900 34804 25956 37212
rect 26012 36372 26068 36382
rect 26012 36370 26292 36372
rect 26012 36318 26014 36370
rect 26066 36318 26292 36370
rect 26012 36316 26292 36318
rect 26012 36306 26068 36316
rect 26236 35810 26292 36316
rect 26236 35758 26238 35810
rect 26290 35758 26292 35810
rect 26236 35746 26292 35758
rect 26796 35700 26852 35710
rect 26796 35606 26852 35644
rect 26908 35308 26964 46508
rect 27804 46562 27972 46564
rect 27804 46510 27918 46562
rect 27970 46510 27972 46562
rect 27804 46508 27972 46510
rect 27804 45892 27860 46508
rect 27916 46498 27972 46508
rect 30716 46564 30772 46622
rect 31500 46676 31556 47182
rect 31500 46620 31780 46676
rect 31164 46564 31220 46574
rect 31276 46564 31332 46574
rect 30716 46562 31332 46564
rect 30716 46510 31166 46562
rect 31218 46510 31278 46562
rect 31330 46510 31332 46562
rect 30716 46508 31332 46510
rect 27020 42868 27076 42878
rect 27020 42082 27076 42812
rect 27020 42030 27022 42082
rect 27074 42030 27076 42082
rect 27020 42018 27076 42030
rect 27468 42532 27524 42542
rect 27468 42084 27524 42476
rect 27468 42018 27524 42028
rect 27804 41860 27860 45836
rect 28812 45220 28868 45230
rect 28812 45126 28868 45164
rect 29036 45106 29092 45118
rect 29036 45054 29038 45106
rect 29090 45054 29092 45106
rect 28140 44996 28196 45006
rect 27916 42756 27972 42766
rect 27916 42662 27972 42700
rect 27468 41804 27860 41860
rect 27020 38834 27076 38846
rect 27020 38782 27022 38834
rect 27074 38782 27076 38834
rect 27020 38612 27076 38782
rect 27468 38834 27524 41804
rect 27468 38782 27470 38834
rect 27522 38782 27524 38834
rect 27468 38770 27524 38782
rect 27692 39620 27748 39630
rect 27692 38668 27748 39564
rect 28140 39618 28196 44940
rect 28476 44996 28532 45006
rect 29036 44996 29092 45054
rect 28476 44994 29092 44996
rect 28476 44942 28478 44994
rect 28530 44942 29092 44994
rect 28476 44940 29092 44942
rect 29260 45108 29316 45118
rect 28364 43652 28420 43662
rect 28364 42980 28420 43596
rect 28364 42754 28420 42924
rect 28364 42702 28366 42754
rect 28418 42702 28420 42754
rect 28364 42690 28420 42702
rect 28140 39566 28142 39618
rect 28194 39566 28196 39618
rect 28140 39554 28196 39566
rect 28364 39620 28420 39630
rect 28364 39526 28420 39564
rect 28476 39396 28532 44940
rect 29260 44322 29316 45052
rect 29596 45108 29652 45118
rect 29596 45014 29652 45052
rect 30716 45108 30772 46508
rect 31164 46470 31220 46508
rect 31276 46498 31332 46508
rect 31724 46562 31780 46620
rect 31724 46510 31726 46562
rect 31778 46510 31780 46562
rect 30716 45042 30772 45052
rect 29260 44270 29262 44322
rect 29314 44270 29316 44322
rect 29260 44258 29316 44270
rect 31612 44994 31668 45006
rect 31612 44942 31614 44994
rect 31666 44942 31668 44994
rect 29932 44210 29988 44222
rect 29932 44158 29934 44210
rect 29986 44158 29988 44210
rect 28812 43652 28868 43662
rect 28812 43558 28868 43596
rect 29260 42756 29316 42766
rect 29260 42662 29316 42700
rect 29484 42754 29540 42766
rect 29484 42702 29486 42754
rect 29538 42702 29540 42754
rect 28588 42532 28644 42542
rect 28588 42438 28644 42476
rect 29484 42532 29540 42702
rect 29708 42756 29764 42766
rect 29708 42662 29764 42700
rect 29484 42466 29540 42476
rect 29596 42532 29652 42542
rect 29932 42532 29988 44158
rect 31500 43428 31556 43438
rect 31612 43428 31668 44942
rect 31500 43426 31668 43428
rect 31500 43374 31502 43426
rect 31554 43374 31668 43426
rect 31500 43372 31668 43374
rect 31500 43316 31556 43372
rect 31500 43250 31556 43260
rect 29596 42530 29988 42532
rect 29596 42478 29598 42530
rect 29650 42478 29988 42530
rect 29596 42476 29988 42478
rect 31388 42980 31444 42990
rect 29596 42466 29652 42476
rect 29820 41972 29876 41982
rect 29148 41860 29204 41870
rect 28924 41804 29148 41860
rect 28140 39340 28532 39396
rect 28588 39506 28644 39518
rect 28588 39454 28590 39506
rect 28642 39454 28644 39506
rect 27020 37828 27076 38556
rect 27020 37762 27076 37772
rect 27132 38612 27748 38668
rect 27916 38722 27972 38734
rect 27916 38670 27918 38722
rect 27970 38670 27972 38722
rect 27132 35924 27188 38612
rect 27916 38388 27972 38670
rect 27916 38322 27972 38332
rect 28140 38050 28196 39340
rect 28476 38722 28532 38734
rect 28476 38670 28478 38722
rect 28530 38670 28532 38722
rect 28476 38612 28532 38670
rect 28476 38546 28532 38556
rect 28588 38276 28644 39454
rect 28588 38210 28644 38220
rect 28140 37998 28142 38050
rect 28194 37998 28196 38050
rect 28140 37986 28196 37998
rect 28364 38050 28420 38062
rect 28364 37998 28366 38050
rect 28418 37998 28420 38050
rect 27244 37826 27300 37838
rect 27244 37774 27246 37826
rect 27298 37774 27300 37826
rect 27244 37716 27300 37774
rect 28364 37716 28420 37998
rect 28588 38052 28644 38062
rect 28588 37958 28644 37996
rect 27244 37660 28420 37716
rect 27132 35858 27188 35868
rect 24668 34354 24724 34748
rect 24668 34302 24670 34354
rect 24722 34302 24724 34354
rect 24668 34290 24724 34302
rect 25228 34802 25620 34804
rect 25228 34750 25342 34802
rect 25394 34750 25620 34802
rect 25228 34748 25620 34750
rect 24332 34244 24388 34254
rect 24332 34150 24388 34188
rect 23772 34018 23828 34030
rect 23772 33966 23774 34018
rect 23826 33966 23828 34018
rect 22540 32732 22932 32788
rect 22652 32564 22708 32574
rect 22092 31106 22204 31108
rect 22092 31054 22094 31106
rect 22146 31054 22204 31106
rect 22092 31052 22204 31054
rect 22092 31042 22148 31052
rect 22204 31014 22260 31052
rect 22540 31106 22596 31118
rect 22540 31054 22542 31106
rect 22594 31054 22596 31106
rect 22316 30996 22372 31006
rect 22316 30902 22372 30940
rect 22540 30884 22596 31054
rect 22652 31106 22708 32508
rect 22652 31054 22654 31106
rect 22706 31054 22708 31106
rect 22652 31042 22708 31054
rect 22764 31220 22820 31230
rect 22540 30818 22596 30828
rect 21980 30382 21982 30434
rect 22034 30382 22036 30434
rect 21980 30370 22036 30382
rect 22204 30380 22708 30436
rect 21756 30146 21812 30156
rect 22092 30212 22148 30222
rect 22204 30212 22260 30380
rect 22092 30210 22260 30212
rect 22092 30158 22094 30210
rect 22146 30158 22260 30210
rect 22092 30156 22260 30158
rect 22316 30212 22372 30222
rect 22092 30146 22148 30156
rect 22316 30118 22372 30156
rect 21532 29988 21588 29998
rect 21980 29988 22036 29998
rect 21532 29986 22036 29988
rect 21532 29934 21534 29986
rect 21586 29934 21982 29986
rect 22034 29934 22036 29986
rect 21532 29932 22036 29934
rect 21532 29922 21588 29932
rect 21980 29876 22036 29932
rect 21980 29810 22036 29820
rect 21420 29596 21812 29652
rect 21756 28084 21812 29596
rect 21308 28082 21812 28084
rect 21308 28030 21758 28082
rect 21810 28030 21812 28082
rect 21308 28028 21812 28030
rect 21308 24948 21364 28028
rect 21756 28018 21812 28028
rect 21868 28532 21924 28542
rect 21868 27970 21924 28476
rect 21868 27918 21870 27970
rect 21922 27918 21924 27970
rect 21868 27906 21924 27918
rect 21532 27858 21588 27870
rect 21532 27806 21534 27858
rect 21586 27806 21588 27858
rect 21420 27076 21476 27086
rect 21532 27076 21588 27806
rect 22428 27860 22484 30380
rect 22652 30210 22708 30380
rect 22652 30158 22654 30210
rect 22706 30158 22708 30210
rect 22652 30146 22708 30158
rect 22540 30100 22596 30110
rect 22540 30006 22596 30044
rect 22652 29652 22708 29662
rect 22652 28756 22708 29596
rect 22540 28532 22596 28542
rect 22540 28438 22596 28476
rect 22652 28530 22708 28700
rect 22652 28478 22654 28530
rect 22706 28478 22708 28530
rect 22652 28466 22708 28478
rect 21980 27636 22036 27646
rect 21420 27074 21588 27076
rect 21420 27022 21422 27074
rect 21474 27022 21588 27074
rect 21420 27020 21588 27022
rect 21644 27074 21700 27086
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 21420 27010 21476 27020
rect 21644 26964 21700 27022
rect 21980 27074 22036 27580
rect 22428 27300 22484 27804
rect 21980 27022 21982 27074
rect 22034 27022 22036 27074
rect 21980 27010 22036 27022
rect 22316 27244 22484 27300
rect 22652 28084 22708 28094
rect 22316 27076 22372 27244
rect 22652 27188 22708 28028
rect 22764 28084 22820 31164
rect 22876 29316 22932 32732
rect 23772 32340 23828 33966
rect 24892 33460 24948 33470
rect 24892 33366 24948 33404
rect 24780 33348 24836 33358
rect 23548 32284 23828 32340
rect 24332 32900 24388 32910
rect 23548 31780 23604 32284
rect 22988 31108 23044 31118
rect 23044 31052 23380 31108
rect 22988 31042 23044 31052
rect 23100 30100 23156 30110
rect 23100 30006 23156 30044
rect 22876 29250 22932 29260
rect 23212 28756 23268 28766
rect 22876 28420 22932 28430
rect 23212 28420 23268 28700
rect 22876 28418 23156 28420
rect 22876 28366 22878 28418
rect 22930 28366 23156 28418
rect 22876 28364 23156 28366
rect 22876 28354 22932 28364
rect 22764 28082 23044 28084
rect 22764 28030 22766 28082
rect 22818 28030 23044 28082
rect 22764 28028 23044 28030
rect 22764 28018 22820 28028
rect 22316 27010 22372 27020
rect 22428 27132 22708 27188
rect 21644 26898 21700 26908
rect 22204 26964 22260 27002
rect 22204 26898 22260 26908
rect 21532 26850 21588 26862
rect 21532 26798 21534 26850
rect 21586 26798 21588 26850
rect 21532 25732 21588 26798
rect 22428 26850 22484 27132
rect 22540 26964 22596 27002
rect 22540 26898 22596 26908
rect 22652 26908 22708 27132
rect 22988 27076 23044 28028
rect 23100 27970 23156 28364
rect 23212 28354 23268 28364
rect 23100 27918 23102 27970
rect 23154 27918 23156 27970
rect 23100 27906 23156 27918
rect 23212 27746 23268 27758
rect 23212 27694 23214 27746
rect 23266 27694 23268 27746
rect 23212 27188 23268 27694
rect 23324 27748 23380 31052
rect 23436 31106 23492 31118
rect 23436 31054 23438 31106
rect 23490 31054 23492 31106
rect 23436 30548 23492 31054
rect 23548 30994 23604 31724
rect 23660 31778 23716 31790
rect 23660 31726 23662 31778
rect 23714 31726 23716 31778
rect 23660 31668 23716 31726
rect 23660 31602 23716 31612
rect 23548 30942 23550 30994
rect 23602 30942 23604 30994
rect 23548 30930 23604 30942
rect 23772 31554 23828 31566
rect 23772 31502 23774 31554
rect 23826 31502 23828 31554
rect 23772 30548 23828 31502
rect 24332 31218 24388 32844
rect 24332 31166 24334 31218
rect 24386 31166 24388 31218
rect 24332 31154 24388 31166
rect 24668 31666 24724 31678
rect 24668 31614 24670 31666
rect 24722 31614 24724 31666
rect 24220 31106 24276 31118
rect 24220 31054 24222 31106
rect 24274 31054 24276 31106
rect 24108 30994 24164 31006
rect 24108 30942 24110 30994
rect 24162 30942 24164 30994
rect 23436 30492 23828 30548
rect 23884 30884 23940 30894
rect 23660 29988 23716 30492
rect 23884 30210 23940 30828
rect 23884 30158 23886 30210
rect 23938 30158 23940 30210
rect 23884 30146 23940 30158
rect 24108 30212 24164 30942
rect 24108 30146 24164 30156
rect 23772 29988 23828 29998
rect 23660 29986 23828 29988
rect 23660 29934 23774 29986
rect 23826 29934 23828 29986
rect 23660 29932 23828 29934
rect 23772 29540 23828 29932
rect 23772 29474 23828 29484
rect 24220 28196 24276 31054
rect 24668 30436 24724 31614
rect 23996 28140 24276 28196
rect 24332 30380 24724 30436
rect 23884 28084 23940 28094
rect 23436 28082 23940 28084
rect 23436 28030 23886 28082
rect 23938 28030 23940 28082
rect 23436 28028 23940 28030
rect 23436 27970 23492 28028
rect 23884 28018 23940 28028
rect 23436 27918 23438 27970
rect 23490 27918 23492 27970
rect 23436 27906 23492 27918
rect 23548 27858 23604 27870
rect 23548 27806 23550 27858
rect 23602 27806 23604 27858
rect 23548 27748 23604 27806
rect 23324 27692 23604 27748
rect 23324 27636 23380 27692
rect 23324 27570 23380 27580
rect 23212 27122 23268 27132
rect 23884 27188 23940 27198
rect 23884 27094 23940 27132
rect 23100 27076 23156 27086
rect 22988 27074 23156 27076
rect 22988 27022 23102 27074
rect 23154 27022 23156 27074
rect 22988 27020 23156 27022
rect 23100 27010 23156 27020
rect 22652 26852 22820 26908
rect 22428 26798 22430 26850
rect 22482 26798 22484 26850
rect 22428 26786 22484 26798
rect 22764 26178 22820 26852
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 21644 25732 21700 25742
rect 21532 25676 21644 25732
rect 21644 25666 21700 25676
rect 22316 25732 22372 25742
rect 21308 24882 21364 24892
rect 22316 24834 22372 25676
rect 22316 24782 22318 24834
rect 22370 24782 22372 24834
rect 22316 24770 22372 24782
rect 22540 24836 22596 24846
rect 22540 24050 22596 24780
rect 22540 23998 22542 24050
rect 22594 23998 22596 24050
rect 22540 23986 22596 23998
rect 21196 23156 21252 23166
rect 21196 23062 21252 23100
rect 21308 21476 21364 21486
rect 21308 21382 21364 21420
rect 21420 19908 21476 19918
rect 21420 19814 21476 19852
rect 22764 17444 22820 26126
rect 22988 24724 23044 24734
rect 22988 24630 23044 24668
rect 23660 24724 23716 24734
rect 23660 24610 23716 24668
rect 23660 24558 23662 24610
rect 23714 24558 23716 24610
rect 23660 22372 23716 24558
rect 23660 22306 23716 22316
rect 23884 21812 23940 21822
rect 23996 21812 24052 28140
rect 24108 27972 24164 27982
rect 24108 27878 24164 27916
rect 24220 27860 24276 27870
rect 24108 26516 24164 26526
rect 24220 26516 24276 27804
rect 24108 26514 24276 26516
rect 24108 26462 24110 26514
rect 24162 26462 24276 26514
rect 24108 26460 24276 26462
rect 24108 26450 24164 26460
rect 24332 22596 24388 30380
rect 24780 30322 24836 33292
rect 25004 31890 25060 31902
rect 25004 31838 25006 31890
rect 25058 31838 25060 31890
rect 24780 30270 24782 30322
rect 24834 30270 24836 30322
rect 24780 30258 24836 30270
rect 24892 31778 24948 31790
rect 24892 31726 24894 31778
rect 24946 31726 24948 31778
rect 24892 30212 24948 31726
rect 25004 31668 25060 31838
rect 25004 31602 25060 31612
rect 25004 30212 25060 30222
rect 24892 30156 25004 30212
rect 25004 30118 25060 30156
rect 24556 30098 24612 30110
rect 24556 30046 24558 30098
rect 24610 30046 24612 30098
rect 24444 26292 24500 26302
rect 24444 26198 24500 26236
rect 23436 21810 24052 21812
rect 23436 21758 23886 21810
rect 23938 21758 24052 21810
rect 23436 21756 24052 21758
rect 24108 22540 24388 22596
rect 23436 21474 23492 21756
rect 23884 21746 23940 21756
rect 23996 21588 24052 21598
rect 23996 21494 24052 21532
rect 23436 21422 23438 21474
rect 23490 21422 23492 21474
rect 23436 21410 23492 21422
rect 23548 21476 23604 21486
rect 23212 20692 23268 20702
rect 22764 17378 22820 17388
rect 23100 20690 23268 20692
rect 23100 20638 23214 20690
rect 23266 20638 23268 20690
rect 23100 20636 23268 20638
rect 23100 19460 23156 20636
rect 23212 20626 23268 20636
rect 23436 20690 23492 20702
rect 23436 20638 23438 20690
rect 23490 20638 23492 20690
rect 23436 19684 23492 20638
rect 23548 20578 23604 21420
rect 23884 21362 23940 21374
rect 24108 21364 24164 22540
rect 24332 22372 24388 22382
rect 23884 21310 23886 21362
rect 23938 21310 23940 21362
rect 23884 20802 23940 21310
rect 23884 20750 23886 20802
rect 23938 20750 23940 20802
rect 23884 20738 23940 20750
rect 23996 21308 24164 21364
rect 24220 21588 24276 21598
rect 23548 20526 23550 20578
rect 23602 20526 23604 20578
rect 23548 20514 23604 20526
rect 23996 20244 24052 21308
rect 23548 20188 24052 20244
rect 23548 19906 23604 20188
rect 23996 20130 24052 20188
rect 23996 20078 23998 20130
rect 24050 20078 24052 20130
rect 23996 20066 24052 20078
rect 24108 20356 24164 20366
rect 24220 20356 24276 21532
rect 24332 21586 24388 22316
rect 24556 21700 24612 30046
rect 24668 28308 24724 28318
rect 24668 28082 24724 28252
rect 24668 28030 24670 28082
rect 24722 28030 24724 28082
rect 24668 27972 24724 28030
rect 24668 23380 24724 27916
rect 24780 24052 24836 24062
rect 24780 23958 24836 23996
rect 24668 23324 24948 23380
rect 24556 21634 24612 21644
rect 24780 23156 24836 23166
rect 24332 21534 24334 21586
rect 24386 21534 24388 21586
rect 24332 21522 24388 21534
rect 24164 20300 24276 20356
rect 24444 21474 24500 21486
rect 24444 21422 24446 21474
rect 24498 21422 24500 21474
rect 24444 21362 24500 21422
rect 24444 21310 24446 21362
rect 24498 21310 24500 21362
rect 23548 19854 23550 19906
rect 23602 19854 23604 19906
rect 23548 19842 23604 19854
rect 23772 20018 23828 20030
rect 23772 19966 23774 20018
rect 23826 19966 23828 20018
rect 23436 19628 23604 19684
rect 23100 19010 23156 19404
rect 23100 18958 23102 19010
rect 23154 18958 23156 19010
rect 21084 16706 21140 16716
rect 21644 16772 21700 16782
rect 21644 16678 21700 16716
rect 23100 16100 23156 18958
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 19012 23380 19182
rect 23324 18946 23380 18956
rect 23436 18004 23492 18014
rect 23100 16006 23156 16044
rect 23324 16772 23380 16782
rect 23212 15986 23268 15998
rect 23212 15934 23214 15986
rect 23266 15934 23268 15986
rect 20972 15250 21028 15260
rect 22092 15316 22148 15326
rect 22092 15222 22148 15260
rect 21644 15202 21700 15214
rect 21644 15150 21646 15202
rect 21698 15150 21700 15202
rect 21644 15148 21700 15150
rect 20972 15092 21700 15148
rect 20972 13858 21028 15092
rect 20972 13806 20974 13858
rect 21026 13806 21028 13858
rect 20972 13794 21028 13806
rect 21756 13636 21812 13646
rect 21756 13542 21812 13580
rect 20860 13524 20916 13534
rect 20860 13430 20916 13468
rect 20412 12014 20414 12066
rect 20466 12014 20468 12066
rect 20412 11508 20468 12014
rect 22876 12740 22932 12750
rect 21420 11508 21476 11518
rect 20412 11506 21476 11508
rect 20412 11454 21422 11506
rect 21474 11454 21476 11506
rect 20412 11452 21476 11454
rect 20412 11394 20468 11452
rect 21420 11442 21476 11452
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20412 11330 20468 11342
rect 20748 11284 20804 11294
rect 20748 11282 20916 11284
rect 20748 11230 20750 11282
rect 20802 11230 20916 11282
rect 20748 11228 20916 11230
rect 20748 11218 20804 11228
rect 19628 11172 19684 11182
rect 19628 10836 19684 11116
rect 20636 11170 20692 11182
rect 20636 11118 20638 11170
rect 20690 11118 20692 11170
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10834 20020 10836
rect 19628 10782 19630 10834
rect 19682 10782 20020 10834
rect 19628 10780 20020 10782
rect 19628 10770 19684 10780
rect 19516 10556 19684 10612
rect 17500 10546 17556 10556
rect 18844 10500 18900 10510
rect 18844 10498 19572 10500
rect 18844 10446 18846 10498
rect 18898 10446 19572 10498
rect 18844 10444 19572 10446
rect 18844 10434 18900 10444
rect 17388 9886 17390 9938
rect 17442 9886 17444 9938
rect 17388 9874 17444 9886
rect 19516 9938 19572 10444
rect 19516 9886 19518 9938
rect 19570 9886 19572 9938
rect 19516 9874 19572 9886
rect 16156 9762 16212 9772
rect 16604 9826 16660 9838
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16268 9604 16324 9614
rect 16604 9604 16660 9774
rect 15708 9602 16660 9604
rect 15708 9550 16270 9602
rect 16322 9550 16660 9602
rect 15708 9548 16660 9550
rect 16716 9604 16772 9614
rect 15372 8370 15540 8372
rect 15372 8318 15374 8370
rect 15426 8318 15540 8370
rect 15372 8316 15540 8318
rect 15372 8306 15428 8316
rect 16268 7364 16324 9548
rect 16716 9266 16772 9548
rect 16716 9214 16718 9266
rect 16770 9214 16772 9266
rect 16716 9202 16772 9214
rect 19628 9156 19684 10556
rect 19964 10610 20020 10780
rect 20636 10724 20692 11118
rect 20748 10724 20804 10734
rect 20636 10722 20804 10724
rect 20636 10670 20750 10722
rect 20802 10670 20804 10722
rect 20636 10668 20804 10670
rect 20748 10658 20804 10668
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19964 10546 20020 10558
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 16828 8932 16884 8942
rect 16828 8930 17556 8932
rect 16828 8878 16830 8930
rect 16882 8878 17556 8930
rect 16828 8876 17556 8878
rect 16828 8866 16884 8876
rect 17500 8370 17556 8876
rect 17500 8318 17502 8370
rect 17554 8318 17556 8370
rect 17500 8306 17556 8318
rect 19628 8260 19684 9100
rect 20860 8596 20916 11228
rect 22876 10500 22932 12684
rect 23212 11618 23268 15934
rect 23324 15874 23380 16716
rect 23324 15822 23326 15874
rect 23378 15822 23380 15874
rect 23324 15810 23380 15822
rect 23436 13412 23492 17948
rect 23548 15148 23604 19628
rect 23772 19234 23828 19966
rect 24108 20018 24164 20300
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 23884 19908 23940 19918
rect 23884 19346 23940 19852
rect 23884 19294 23886 19346
rect 23938 19294 23940 19346
rect 23884 19282 23940 19294
rect 24108 19348 24164 19966
rect 24444 19908 24500 21310
rect 24780 20020 24836 23100
rect 24556 19908 24612 19918
rect 24444 19906 24612 19908
rect 24444 19854 24558 19906
rect 24610 19854 24612 19906
rect 24444 19852 24612 19854
rect 24108 19282 24164 19292
rect 24444 19348 24500 19358
rect 23772 19182 23774 19234
rect 23826 19182 23828 19234
rect 23772 19170 23828 19182
rect 23996 19236 24052 19246
rect 23996 19142 24052 19180
rect 24332 19122 24388 19134
rect 24332 19070 24334 19122
rect 24386 19070 24388 19122
rect 24332 19012 24388 19070
rect 24332 18946 24388 18956
rect 24332 17556 24388 17566
rect 23772 17108 23828 17118
rect 23772 16770 23828 17052
rect 24220 17108 24276 17118
rect 24220 17014 24276 17052
rect 24332 16994 24388 17500
rect 24332 16942 24334 16994
rect 24386 16942 24388 16994
rect 24332 16930 24388 16942
rect 23996 16884 24052 16894
rect 23772 16718 23774 16770
rect 23826 16718 23828 16770
rect 23772 16706 23828 16718
rect 23884 16882 24052 16884
rect 23884 16830 23998 16882
rect 24050 16830 24052 16882
rect 23884 16828 24052 16830
rect 23884 16324 23940 16828
rect 23996 16818 24052 16828
rect 23660 16268 23940 16324
rect 24108 16772 24164 16782
rect 23660 16098 23716 16268
rect 23660 16046 23662 16098
rect 23714 16046 23716 16098
rect 23660 16034 23716 16046
rect 23996 15876 24052 15886
rect 24108 15876 24164 16716
rect 24444 16098 24500 19292
rect 24556 19236 24612 19852
rect 24556 19170 24612 19180
rect 24780 19012 24836 19964
rect 24556 19010 24836 19012
rect 24556 18958 24782 19010
rect 24834 18958 24836 19010
rect 24556 18956 24836 18958
rect 24556 18674 24612 18956
rect 24780 18946 24836 18956
rect 24556 18622 24558 18674
rect 24610 18622 24612 18674
rect 24556 18610 24612 18622
rect 24892 18340 24948 23324
rect 25004 22260 25060 22270
rect 25004 22166 25060 22204
rect 25228 20916 25284 34748
rect 25340 34738 25396 34748
rect 25564 34580 25620 34748
rect 25732 34748 25956 34804
rect 26572 35252 26964 35308
rect 27132 35586 27188 35598
rect 27132 35534 27134 35586
rect 27186 35534 27188 35586
rect 27132 35364 27188 35534
rect 27132 35298 27188 35308
rect 25676 34710 25732 34748
rect 26124 34690 26180 34702
rect 26124 34638 26126 34690
rect 26178 34638 26180 34690
rect 26124 34580 26180 34638
rect 25564 34524 26180 34580
rect 25564 33460 25620 33470
rect 25564 32786 25620 33404
rect 25564 32734 25566 32786
rect 25618 32734 25620 32786
rect 25452 32564 25508 32574
rect 25340 32508 25452 32564
rect 25340 30098 25396 32508
rect 25452 32470 25508 32508
rect 25564 32452 25620 32734
rect 26236 33236 26292 33246
rect 26236 32786 26292 33180
rect 26236 32734 26238 32786
rect 26290 32734 26292 32786
rect 26236 32722 26292 32734
rect 25788 32674 25844 32686
rect 25788 32622 25790 32674
rect 25842 32622 25844 32674
rect 25788 32564 25844 32622
rect 25900 32564 25956 32574
rect 25788 32562 25956 32564
rect 25788 32510 25902 32562
rect 25954 32510 25956 32562
rect 25788 32508 25956 32510
rect 25900 32498 25956 32508
rect 26236 32562 26292 32574
rect 26236 32510 26238 32562
rect 26290 32510 26292 32562
rect 25564 32386 25620 32396
rect 26012 31556 26068 31566
rect 25340 30046 25342 30098
rect 25394 30046 25396 30098
rect 25340 30034 25396 30046
rect 25452 31108 25508 31118
rect 25452 30100 25508 31052
rect 26012 30324 26068 31500
rect 26012 30258 26068 30268
rect 26124 30212 26180 30222
rect 26236 30212 26292 32510
rect 26348 32564 26404 32574
rect 26348 31778 26404 32508
rect 26572 32562 26628 35252
rect 27132 34130 27188 34142
rect 27132 34078 27134 34130
rect 27186 34078 27188 34130
rect 27132 34020 27188 34078
rect 27804 34020 27860 34030
rect 27132 33954 27188 33964
rect 27244 34018 27860 34020
rect 27244 33966 27806 34018
rect 27858 33966 27860 34018
rect 27244 33964 27860 33966
rect 27020 33236 27076 33246
rect 27020 33142 27076 33180
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 26572 32452 26628 32510
rect 27020 32452 27076 32462
rect 26572 32450 27076 32452
rect 26572 32398 27022 32450
rect 27074 32398 27076 32450
rect 26572 32396 27076 32398
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26348 31714 26404 31726
rect 26684 31780 26740 31790
rect 26908 31780 26964 31790
rect 26684 31778 26964 31780
rect 26684 31726 26686 31778
rect 26738 31726 26910 31778
rect 26962 31726 26964 31778
rect 26684 31724 26964 31726
rect 26684 31714 26740 31724
rect 26908 31714 26964 31724
rect 26460 31556 26516 31566
rect 26460 31462 26516 31500
rect 26684 31332 26740 31342
rect 26684 31218 26740 31276
rect 27020 31332 27076 32396
rect 27244 31554 27300 33964
rect 27804 33954 27860 33964
rect 28252 34020 28308 34030
rect 28252 33460 28308 33964
rect 27804 33458 28308 33460
rect 27804 33406 28254 33458
rect 28306 33406 28308 33458
rect 27804 33404 28308 33406
rect 27804 33346 27860 33404
rect 28252 33394 28308 33404
rect 27804 33294 27806 33346
rect 27858 33294 27860 33346
rect 27804 33282 27860 33294
rect 28364 33236 28420 37660
rect 28812 37268 28868 37278
rect 28924 37268 28980 41804
rect 29148 41766 29204 41804
rect 29372 41860 29428 41870
rect 29260 39620 29316 39630
rect 29260 39394 29316 39564
rect 29260 39342 29262 39394
rect 29314 39342 29316 39394
rect 29148 38946 29204 38958
rect 29148 38894 29150 38946
rect 29202 38894 29204 38946
rect 29036 38834 29092 38846
rect 29036 38782 29038 38834
rect 29090 38782 29092 38834
rect 29036 37492 29092 38782
rect 29148 38274 29204 38894
rect 29260 38836 29316 39342
rect 29372 39058 29428 41804
rect 29372 39006 29374 39058
rect 29426 39006 29428 39058
rect 29372 38994 29428 39006
rect 29820 40404 29876 41916
rect 30380 41972 30436 41982
rect 30380 41186 30436 41916
rect 30380 41134 30382 41186
rect 30434 41134 30436 41186
rect 30380 41122 30436 41134
rect 31052 41076 31108 41086
rect 31052 40982 31108 41020
rect 30044 40628 30100 40638
rect 30380 40628 30436 40638
rect 30100 40626 30436 40628
rect 30100 40574 30382 40626
rect 30434 40574 30436 40626
rect 30100 40572 30436 40574
rect 30044 40534 30100 40572
rect 30380 40562 30436 40572
rect 30716 40628 30772 40638
rect 30716 40534 30772 40572
rect 31388 40626 31444 42924
rect 31724 42980 31780 46510
rect 31836 46452 31892 46462
rect 31948 46452 32004 47292
rect 32620 47348 32676 47358
rect 32620 47346 33124 47348
rect 32620 47294 32622 47346
rect 32674 47294 33124 47346
rect 32620 47292 33124 47294
rect 32620 47282 32676 47292
rect 33068 46562 33124 47292
rect 33180 47236 33236 47246
rect 33180 46898 33236 47180
rect 33180 46846 33182 46898
rect 33234 46846 33236 46898
rect 33180 46834 33236 46846
rect 33404 46786 33460 48076
rect 33404 46734 33406 46786
rect 33458 46734 33460 46786
rect 33404 46722 33460 46734
rect 33068 46510 33070 46562
rect 33122 46510 33124 46562
rect 33068 46498 33124 46510
rect 31836 46450 32228 46452
rect 31836 46398 31838 46450
rect 31890 46398 32228 46450
rect 31836 46396 32228 46398
rect 31836 46386 31892 46396
rect 31724 42914 31780 42924
rect 31948 45106 32004 45118
rect 31948 45054 31950 45106
rect 32002 45054 32004 45106
rect 31948 44436 32004 45054
rect 31948 43314 32004 44380
rect 32060 44548 32116 44558
rect 32060 44434 32116 44492
rect 32060 44382 32062 44434
rect 32114 44382 32116 44434
rect 32060 44370 32116 44382
rect 32172 43428 32228 46396
rect 33068 45220 33124 45230
rect 33068 45126 33124 45164
rect 32396 45108 32452 45118
rect 32396 45014 32452 45052
rect 33628 45106 33684 45118
rect 33628 45054 33630 45106
rect 33682 45054 33684 45106
rect 33516 44884 33572 44894
rect 33404 44828 33516 44884
rect 33292 44548 33348 44558
rect 33404 44548 33460 44828
rect 33516 44818 33572 44828
rect 33628 44548 33684 45054
rect 33852 45108 33908 45118
rect 33852 44994 33908 45052
rect 33852 44942 33854 44994
rect 33906 44942 33908 44994
rect 33852 44930 33908 44942
rect 33292 44546 33460 44548
rect 33292 44494 33294 44546
rect 33346 44494 33460 44546
rect 33292 44492 33460 44494
rect 33516 44492 33684 44548
rect 33852 44548 33908 44558
rect 33292 44482 33348 44492
rect 32732 44436 32788 44446
rect 32788 44380 32900 44436
rect 32732 44370 32788 44380
rect 32396 44324 32452 44334
rect 32284 44268 32396 44324
rect 32284 43538 32340 44268
rect 32396 44230 32452 44268
rect 32620 44322 32676 44334
rect 32620 44270 32622 44322
rect 32674 44270 32676 44322
rect 32284 43486 32286 43538
rect 32338 43486 32340 43538
rect 32284 43474 32340 43486
rect 31948 43262 31950 43314
rect 32002 43262 32004 43314
rect 31948 41860 32004 43262
rect 32060 43316 32116 43326
rect 32060 42868 32116 43260
rect 32172 43092 32228 43372
rect 32396 43426 32452 43438
rect 32396 43374 32398 43426
rect 32450 43374 32452 43426
rect 32396 43316 32452 43374
rect 32396 43250 32452 43260
rect 32172 43036 32452 43092
rect 32060 42802 32116 42812
rect 32396 42866 32452 43036
rect 32396 42814 32398 42866
rect 32450 42814 32452 42866
rect 32396 42802 32452 42814
rect 32620 42868 32676 44270
rect 32844 44322 32900 44380
rect 32844 44270 32846 44322
rect 32898 44270 32900 44322
rect 32844 44258 32900 44270
rect 33516 44212 33572 44492
rect 33628 44324 33684 44334
rect 33684 44268 33796 44324
rect 33628 44230 33684 44268
rect 33068 43538 33124 43550
rect 33068 43486 33070 43538
rect 33122 43486 33124 43538
rect 32732 42868 32788 42878
rect 33068 42868 33124 43486
rect 33516 43426 33572 44156
rect 33516 43374 33518 43426
rect 33570 43374 33572 43426
rect 33516 43362 33572 43374
rect 33740 42978 33796 44268
rect 33740 42926 33742 42978
rect 33794 42926 33796 42978
rect 33740 42914 33796 42926
rect 32620 42812 32732 42868
rect 32788 42812 33124 42868
rect 33852 42866 33908 44492
rect 33964 42980 34020 48748
rect 34300 48244 34356 49420
rect 34524 48468 34580 48478
rect 34748 48468 34804 49756
rect 34524 48466 34804 48468
rect 34524 48414 34526 48466
rect 34578 48414 34804 48466
rect 34524 48412 34804 48414
rect 34860 49810 34916 49822
rect 34860 49758 34862 49810
rect 34914 49758 34916 49810
rect 34860 48692 34916 49758
rect 35084 49810 35140 49980
rect 36764 50036 36820 50372
rect 36764 49942 36820 49980
rect 37212 50036 37268 50046
rect 37212 49922 37268 49980
rect 37660 50034 37716 50428
rect 39116 50484 39172 50494
rect 39116 50390 39172 50428
rect 37660 49982 37662 50034
rect 37714 49982 37716 50034
rect 37660 49970 37716 49982
rect 39788 50036 39844 50046
rect 40236 50036 40292 50654
rect 39844 49980 40292 50036
rect 41020 50484 41076 50494
rect 41020 50034 41076 50428
rect 41020 49982 41022 50034
rect 41074 49982 41076 50034
rect 37212 49870 37214 49922
rect 37266 49870 37268 49922
rect 37212 49858 37268 49870
rect 37772 49924 37828 49934
rect 37772 49830 37828 49868
rect 35084 49758 35086 49810
rect 35138 49758 35140 49810
rect 35084 48804 35140 49758
rect 36652 49812 36708 49822
rect 36652 49718 36708 49756
rect 36988 49810 37044 49822
rect 36988 49758 36990 49810
rect 37042 49758 37044 49810
rect 36876 49700 36932 49710
rect 36876 49606 36932 49644
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35084 48738 35140 48748
rect 34860 48466 34916 48636
rect 34860 48414 34862 48466
rect 34914 48414 34916 48466
rect 34524 48402 34580 48412
rect 34860 48402 34916 48414
rect 36988 48692 37044 49758
rect 39004 49812 39060 49822
rect 39564 49812 39620 49822
rect 39060 49810 39620 49812
rect 39060 49758 39566 49810
rect 39618 49758 39620 49810
rect 39060 49756 39620 49758
rect 37548 49700 37604 49710
rect 37548 49606 37604 49644
rect 37772 48916 37828 48926
rect 37828 48860 37940 48916
rect 37772 48850 37828 48860
rect 34188 45106 34244 45118
rect 34188 45054 34190 45106
rect 34242 45054 34244 45106
rect 34188 44548 34244 45054
rect 34188 44482 34244 44492
rect 34076 44324 34132 44334
rect 34076 44322 34244 44324
rect 34076 44270 34078 44322
rect 34130 44270 34244 44322
rect 34076 44268 34244 44270
rect 34076 44258 34132 44268
rect 34188 43876 34244 44268
rect 34188 43538 34244 43820
rect 34188 43486 34190 43538
rect 34242 43486 34244 43538
rect 34188 43474 34244 43486
rect 34188 43314 34244 43326
rect 34188 43262 34190 43314
rect 34242 43262 34244 43314
rect 34188 43204 34244 43262
rect 34188 43138 34244 43148
rect 34076 42980 34132 42990
rect 33964 42978 34132 42980
rect 33964 42926 34078 42978
rect 34130 42926 34132 42978
rect 33964 42924 34132 42926
rect 34076 42914 34132 42924
rect 33852 42814 33854 42866
rect 33906 42814 33908 42866
rect 32732 42774 32788 42812
rect 33852 42802 33908 42814
rect 33628 42532 33684 42542
rect 33628 42308 33684 42476
rect 33404 42252 33684 42308
rect 33404 42082 33460 42252
rect 33404 42030 33406 42082
rect 33458 42030 33460 42082
rect 33404 42018 33460 42030
rect 33516 42082 33572 42094
rect 33516 42030 33518 42082
rect 33570 42030 33572 42082
rect 31948 41794 32004 41804
rect 33180 41300 33236 41310
rect 33516 41300 33572 42030
rect 31388 40574 31390 40626
rect 31442 40574 31444 40626
rect 31388 40562 31444 40574
rect 33068 41298 33572 41300
rect 33068 41246 33182 41298
rect 33234 41246 33572 41298
rect 33068 41244 33572 41246
rect 33628 41300 33684 42252
rect 34300 42196 34356 48188
rect 34636 48244 34692 48254
rect 34972 48244 35028 48254
rect 34636 48242 34804 48244
rect 34636 48190 34638 48242
rect 34690 48190 34804 48242
rect 34636 48188 34804 48190
rect 34636 48178 34692 48188
rect 34524 48132 34580 48142
rect 34524 48038 34580 48076
rect 34748 47570 34804 48188
rect 34972 48150 35028 48188
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34748 47518 34750 47570
rect 34802 47518 34804 47570
rect 34748 47068 34804 47518
rect 35196 47348 35252 47358
rect 35196 47254 35252 47292
rect 36988 47346 37044 48636
rect 37772 47684 37828 47694
rect 37772 47590 37828 47628
rect 36988 47294 36990 47346
rect 37042 47294 37044 47346
rect 34748 47012 35028 47068
rect 34748 46004 34804 46014
rect 34524 46002 34804 46004
rect 34524 45950 34750 46002
rect 34802 45950 34804 46002
rect 34524 45948 34804 45950
rect 34412 44210 34468 44222
rect 34412 44158 34414 44210
rect 34466 44158 34468 44210
rect 34412 43652 34468 44158
rect 34412 43586 34468 43596
rect 34524 43650 34580 45948
rect 34748 45938 34804 45948
rect 34860 45668 34916 45678
rect 34636 45666 34916 45668
rect 34636 45614 34862 45666
rect 34914 45614 34916 45666
rect 34636 45612 34916 45614
rect 34636 44212 34692 45612
rect 34860 45602 34916 45612
rect 34860 44996 34916 45006
rect 34748 44548 34804 44558
rect 34748 44322 34804 44492
rect 34748 44270 34750 44322
rect 34802 44270 34804 44322
rect 34748 44258 34804 44270
rect 34636 44146 34692 44156
rect 34524 43598 34526 43650
rect 34578 43598 34580 43650
rect 34524 43586 34580 43598
rect 34860 43540 34916 44940
rect 34748 43538 34916 43540
rect 34748 43486 34862 43538
rect 34914 43486 34916 43538
rect 34748 43484 34916 43486
rect 34524 42756 34580 42766
rect 34412 42532 34468 42542
rect 34412 42438 34468 42476
rect 34412 42196 34468 42206
rect 34300 42194 34468 42196
rect 34300 42142 34414 42194
rect 34466 42142 34468 42194
rect 34300 42140 34468 42142
rect 34412 42130 34468 42140
rect 34524 42084 34580 42700
rect 34524 41990 34580 42028
rect 34748 42530 34804 43484
rect 34860 43474 34916 43484
rect 34748 42478 34750 42530
rect 34802 42478 34804 42530
rect 30604 40516 30660 40526
rect 29708 38836 29764 38846
rect 29820 38836 29876 40348
rect 30492 40460 30604 40516
rect 30380 38948 30436 38958
rect 30492 38948 30548 40460
rect 30604 40450 30660 40460
rect 31052 40402 31108 40414
rect 31052 40350 31054 40402
rect 31106 40350 31108 40402
rect 30716 39396 30772 39406
rect 31052 39396 31108 40350
rect 30716 39394 31108 39396
rect 30716 39342 30718 39394
rect 30770 39342 31108 39394
rect 30716 39340 31108 39342
rect 32508 39396 32564 39406
rect 30716 39060 30772 39340
rect 30716 38994 30772 39004
rect 30380 38946 30548 38948
rect 30380 38894 30382 38946
rect 30434 38894 30548 38946
rect 30380 38892 30548 38894
rect 30380 38882 30436 38892
rect 29260 38780 29428 38836
rect 29372 38724 29428 38780
rect 29708 38834 29876 38836
rect 29708 38782 29710 38834
rect 29762 38782 29876 38834
rect 29708 38780 29876 38782
rect 29708 38770 29764 38780
rect 32508 38722 32564 39340
rect 32508 38670 32510 38722
rect 32562 38670 32564 38722
rect 32508 38668 32564 38670
rect 33068 38668 33124 41244
rect 33180 41234 33236 41244
rect 29372 38658 29428 38668
rect 32172 38612 32564 38668
rect 32956 38612 33124 38668
rect 33180 40404 33236 40414
rect 33180 40292 33236 40348
rect 33404 40292 33460 40302
rect 33180 40290 33460 40292
rect 33180 40238 33406 40290
rect 33458 40238 33460 40290
rect 33180 40236 33460 40238
rect 33180 39058 33236 40236
rect 33404 40226 33460 40236
rect 33516 39620 33572 39630
rect 33628 39620 33684 41244
rect 33740 41970 33796 41982
rect 33740 41918 33742 41970
rect 33794 41918 33796 41970
rect 33740 41186 33796 41918
rect 34188 41970 34244 41982
rect 34188 41918 34190 41970
rect 34242 41918 34244 41970
rect 33740 41134 33742 41186
rect 33794 41134 33796 41186
rect 33740 41122 33796 41134
rect 34076 41748 34132 41758
rect 34076 41186 34132 41692
rect 34076 41134 34078 41186
rect 34130 41134 34132 41186
rect 34076 41122 34132 41134
rect 33852 41076 33908 41086
rect 33852 40982 33908 41020
rect 33964 40516 34020 40526
rect 33964 40422 34020 40460
rect 34188 40514 34244 41918
rect 34188 40462 34190 40514
rect 34242 40462 34244 40514
rect 34188 40450 34244 40462
rect 34300 41076 34356 41086
rect 34300 40628 34356 41020
rect 33572 39564 33684 39620
rect 33852 40402 33908 40414
rect 33852 40350 33854 40402
rect 33906 40350 33908 40402
rect 33852 39618 33908 40350
rect 34300 40402 34356 40572
rect 34300 40350 34302 40402
rect 34354 40350 34356 40402
rect 34300 40338 34356 40350
rect 33852 39566 33854 39618
rect 33906 39566 33908 39618
rect 33516 39526 33572 39564
rect 33852 39554 33908 39566
rect 34188 39620 34244 39630
rect 34188 39526 34244 39564
rect 33628 39396 33684 39406
rect 33628 39302 33684 39340
rect 33180 39006 33182 39058
rect 33234 39006 33236 39058
rect 29820 38388 29876 38398
rect 29148 38222 29150 38274
rect 29202 38222 29204 38274
rect 29148 38210 29204 38222
rect 29708 38276 29764 38286
rect 29708 38182 29764 38220
rect 29820 38274 29876 38332
rect 29820 38222 29822 38274
rect 29874 38222 29876 38274
rect 29820 38210 29876 38222
rect 29036 37426 29092 37436
rect 29260 38050 29316 38062
rect 29260 37998 29262 38050
rect 29314 37998 29316 38050
rect 29260 37378 29316 37998
rect 29484 38052 29540 38062
rect 29484 37958 29540 37996
rect 29260 37326 29262 37378
rect 29314 37326 29316 37378
rect 29260 37314 29316 37326
rect 30828 37380 30884 37390
rect 28812 37266 28980 37268
rect 28812 37214 28814 37266
rect 28866 37214 28980 37266
rect 28812 37212 28980 37214
rect 29148 37266 29204 37278
rect 29148 37214 29150 37266
rect 29202 37214 29204 37266
rect 28812 37202 28868 37212
rect 29148 37156 29204 37214
rect 29820 37156 29876 37166
rect 29148 37154 29876 37156
rect 29148 37102 29822 37154
rect 29874 37102 29876 37154
rect 29148 37100 29876 37102
rect 29820 36260 29876 37100
rect 30156 36260 30212 36270
rect 29820 36204 30156 36260
rect 29036 35586 29092 35598
rect 29036 35534 29038 35586
rect 29090 35534 29092 35586
rect 29036 34804 29092 35534
rect 29484 35588 29540 35598
rect 29484 35494 29540 35532
rect 29036 34738 29092 34748
rect 29484 35028 29540 35038
rect 28252 33180 28420 33236
rect 29484 33458 29540 34972
rect 29484 33406 29486 33458
rect 29538 33406 29540 33458
rect 27916 32452 27972 32462
rect 27468 31778 27524 31790
rect 27468 31726 27470 31778
rect 27522 31726 27524 31778
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 27244 31490 27300 31502
rect 27356 31666 27412 31678
rect 27356 31614 27358 31666
rect 27410 31614 27412 31666
rect 27020 31266 27076 31276
rect 26684 31166 26686 31218
rect 26738 31166 26740 31218
rect 26684 31154 26740 31166
rect 27356 31218 27412 31614
rect 27356 31166 27358 31218
rect 27410 31166 27412 31218
rect 27356 31154 27412 31166
rect 27468 31332 27524 31726
rect 27916 31778 27972 32396
rect 27916 31726 27918 31778
rect 27970 31726 27972 31778
rect 27916 31714 27972 31726
rect 28140 31556 28196 31566
rect 28140 31462 28196 31500
rect 26124 30210 26292 30212
rect 26124 30158 26126 30210
rect 26178 30158 26292 30210
rect 26124 30156 26292 30158
rect 26460 30996 26516 31006
rect 26124 30146 26180 30156
rect 25452 30034 25508 30044
rect 26460 30098 26516 30940
rect 26460 30046 26462 30098
rect 26514 30046 26516 30098
rect 25676 29986 25732 29998
rect 25676 29934 25678 29986
rect 25730 29934 25732 29986
rect 25676 28532 25732 29934
rect 26348 29988 26404 29998
rect 26348 29894 26404 29932
rect 26460 29540 26516 30046
rect 27020 29988 27076 29998
rect 27020 29894 27076 29932
rect 25676 27300 25732 28476
rect 26348 29484 26516 29540
rect 26908 29650 26964 29662
rect 26908 29598 26910 29650
rect 26962 29598 26964 29650
rect 26908 29540 26964 29598
rect 26964 29484 27076 29540
rect 25676 27234 25732 27244
rect 26012 28420 26068 28430
rect 26012 27186 26068 28364
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27122 26068 27134
rect 26348 26908 26404 29484
rect 26908 29474 26964 29484
rect 26796 29426 26852 29438
rect 26796 29374 26798 29426
rect 26850 29374 26852 29426
rect 26460 29316 26516 29326
rect 26796 29316 26852 29374
rect 26460 29314 26852 29316
rect 26460 29262 26462 29314
rect 26514 29262 26852 29314
rect 26460 29260 26852 29262
rect 26460 28420 26516 29260
rect 27020 28754 27076 29484
rect 27020 28702 27022 28754
rect 27074 28702 27076 28754
rect 27020 28690 27076 28702
rect 27132 28868 27188 28878
rect 26460 28354 26516 28364
rect 26236 26852 26404 26908
rect 26796 28196 26852 28206
rect 25900 26292 25956 26302
rect 25900 25508 25956 26236
rect 25900 25414 25956 25452
rect 26236 25396 26292 26852
rect 26796 26514 26852 28140
rect 26908 27748 26964 27758
rect 26908 27654 26964 27692
rect 27132 26908 27188 28812
rect 27244 27858 27300 27870
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 27244 27748 27300 27806
rect 27244 27682 27300 27692
rect 26796 26462 26798 26514
rect 26850 26462 26852 26514
rect 26796 26450 26852 26462
rect 26908 26852 27188 26908
rect 26908 26292 26964 26852
rect 27468 26516 27524 31276
rect 27580 31106 27636 31118
rect 27580 31054 27582 31106
rect 27634 31054 27636 31106
rect 27580 30884 27636 31054
rect 27692 30996 27748 31006
rect 27692 30902 27748 30940
rect 28140 30996 28196 31006
rect 28140 30902 28196 30940
rect 27580 30818 27636 30828
rect 28252 30772 28308 33180
rect 28588 32116 28644 32126
rect 28588 32004 28644 32060
rect 28476 31948 28644 32004
rect 28476 31890 28532 31948
rect 28476 31838 28478 31890
rect 28530 31838 28532 31890
rect 28476 31826 28532 31838
rect 28588 31780 28644 31790
rect 29484 31780 29540 33406
rect 28588 31778 28756 31780
rect 28588 31726 28590 31778
rect 28642 31726 28756 31778
rect 28588 31724 28756 31726
rect 28588 31714 28644 31724
rect 28140 30716 28308 30772
rect 28364 31554 28420 31566
rect 28364 31502 28366 31554
rect 28418 31502 28420 31554
rect 28028 29986 28084 29998
rect 28028 29934 28030 29986
rect 28082 29934 28084 29986
rect 27916 29652 27972 29662
rect 27916 29558 27972 29596
rect 27804 29538 27860 29550
rect 27804 29486 27806 29538
rect 27858 29486 27860 29538
rect 27580 28644 27636 28654
rect 27580 28550 27636 28588
rect 27580 27300 27636 27310
rect 27580 27206 27636 27244
rect 27692 26962 27748 26974
rect 27692 26910 27694 26962
rect 27746 26910 27748 26962
rect 27580 26852 27636 26862
rect 27580 26758 27636 26796
rect 27692 26740 27748 26910
rect 27692 26674 27748 26684
rect 27580 26516 27636 26526
rect 27468 26460 27580 26516
rect 27580 26450 27636 26460
rect 27804 26292 27860 29486
rect 28028 29316 28084 29934
rect 28028 28644 28084 29260
rect 28140 28868 28196 30716
rect 28140 28802 28196 28812
rect 28252 29426 28308 29438
rect 28252 29374 28254 29426
rect 28306 29374 28308 29426
rect 27916 28420 27972 28430
rect 27916 28196 27972 28364
rect 27916 28130 27972 28140
rect 28028 28418 28084 28588
rect 28028 28366 28030 28418
rect 28082 28366 28084 28418
rect 28028 26908 28084 28366
rect 28252 28196 28308 29374
rect 28252 28130 28308 28140
rect 28364 26908 28420 31502
rect 28588 31556 28644 31566
rect 28588 30322 28644 31500
rect 28588 30270 28590 30322
rect 28642 30270 28644 30322
rect 28588 30258 28644 30270
rect 28700 30212 28756 31724
rect 29484 31714 29540 31724
rect 29708 34804 29764 34814
rect 29708 34690 29764 34748
rect 29708 34638 29710 34690
rect 29762 34638 29764 34690
rect 29260 31556 29316 31566
rect 29260 31462 29316 31500
rect 29708 31556 29764 34638
rect 29708 31490 29764 31500
rect 29932 34692 29988 34702
rect 29932 34018 29988 34636
rect 29932 33966 29934 34018
rect 29986 33966 29988 34018
rect 29596 31332 29652 31342
rect 28700 30146 28756 30156
rect 29148 30212 29204 30222
rect 29148 30118 29204 30156
rect 29596 29652 29652 31276
rect 29932 31220 29988 33966
rect 29932 31154 29988 31164
rect 29708 30100 29764 30110
rect 29708 30006 29764 30044
rect 29596 29586 29652 29596
rect 28812 29316 28868 29326
rect 28812 29222 28868 29260
rect 28028 26852 28196 26908
rect 28140 26850 28196 26852
rect 28140 26798 28142 26850
rect 28194 26798 28196 26850
rect 28140 26740 28196 26798
rect 26684 26236 26964 26292
rect 27244 26236 27860 26292
rect 28028 26516 28084 26526
rect 26124 25394 26292 25396
rect 26124 25342 26238 25394
rect 26290 25342 26292 25394
rect 26124 25340 26292 25342
rect 25564 25284 25620 25294
rect 25564 24836 25620 25228
rect 25564 24770 25620 24780
rect 26124 24836 26180 25340
rect 26236 25330 26292 25340
rect 26572 25508 26628 25518
rect 26684 25508 26740 26236
rect 26572 25506 26740 25508
rect 26572 25454 26574 25506
rect 26626 25454 26740 25506
rect 26572 25452 26740 25454
rect 27132 25732 27188 25742
rect 26572 25284 26628 25452
rect 26908 25394 26964 25406
rect 26908 25342 26910 25394
rect 26962 25342 26964 25394
rect 26572 25218 26628 25228
rect 26796 25282 26852 25294
rect 26796 25230 26798 25282
rect 26850 25230 26852 25282
rect 26124 24742 26180 24780
rect 26460 25172 26516 25182
rect 26460 24722 26516 25116
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 26460 24658 26516 24670
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24052 26292 24558
rect 26684 24500 26740 24510
rect 26796 24500 26852 25230
rect 26908 25284 26964 25342
rect 26908 25218 26964 25228
rect 27132 25172 27188 25676
rect 26684 24498 26852 24500
rect 26684 24446 26686 24498
rect 26738 24446 26852 24498
rect 26684 24444 26852 24446
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26908 24612 26964 24670
rect 26684 24434 26740 24444
rect 26236 23986 26292 23996
rect 25564 23938 25620 23950
rect 25564 23886 25566 23938
rect 25618 23886 25620 23938
rect 25564 23716 25620 23886
rect 26908 23828 26964 24556
rect 27132 24050 27188 25116
rect 27132 23998 27134 24050
rect 27186 23998 27188 24050
rect 27132 23986 27188 23998
rect 26684 23772 26964 23828
rect 26012 23716 26068 23726
rect 25564 23714 26068 23716
rect 25564 23662 26014 23714
rect 26066 23662 26068 23714
rect 25564 23660 26068 23662
rect 26012 23044 26068 23660
rect 26012 22372 26068 22988
rect 26012 22306 26068 22316
rect 25228 20850 25284 20860
rect 26684 20132 26740 23772
rect 27132 22484 27188 22494
rect 27244 22484 27300 26236
rect 27692 25508 27748 25518
rect 27916 25508 27972 25518
rect 27692 25506 27916 25508
rect 27692 25454 27694 25506
rect 27746 25454 27916 25506
rect 27692 25452 27916 25454
rect 27692 25442 27748 25452
rect 27916 25414 27972 25452
rect 27468 24612 27524 24622
rect 27468 24518 27524 24556
rect 27356 23044 27412 23054
rect 27356 22950 27412 22988
rect 26908 22482 27300 22484
rect 26908 22430 27134 22482
rect 27186 22430 27300 22482
rect 26908 22428 27300 22430
rect 26908 21810 26964 22428
rect 27132 22418 27188 22428
rect 27356 22372 27412 22382
rect 27244 22370 27412 22372
rect 27244 22318 27358 22370
rect 27410 22318 27412 22370
rect 27244 22316 27412 22318
rect 26908 21758 26910 21810
rect 26962 21758 26964 21810
rect 26908 21746 26964 21758
rect 27132 21812 27188 21822
rect 27244 21812 27300 22316
rect 27356 22306 27412 22316
rect 27692 22370 27748 22382
rect 28028 22372 28084 26460
rect 28140 25506 28196 26684
rect 28140 25454 28142 25506
rect 28194 25454 28196 25506
rect 28140 25396 28196 25454
rect 28140 25330 28196 25340
rect 28252 26852 28420 26908
rect 28588 28532 28644 28542
rect 28140 24612 28196 24622
rect 28140 24518 28196 24556
rect 27692 22318 27694 22370
rect 27746 22318 27748 22370
rect 27580 22260 27636 22270
rect 27580 22166 27636 22204
rect 27692 22036 27748 22318
rect 27132 21810 27300 21812
rect 27132 21758 27134 21810
rect 27186 21758 27300 21810
rect 27132 21756 27300 21758
rect 27468 21980 27748 22036
rect 27804 22370 28084 22372
rect 27804 22318 28030 22370
rect 28082 22318 28084 22370
rect 27804 22316 28084 22318
rect 27132 21746 27188 21756
rect 26796 21586 26852 21598
rect 26796 21534 26798 21586
rect 26850 21534 26852 21586
rect 26796 20356 26852 21534
rect 26796 20290 26852 20300
rect 26796 20132 26852 20142
rect 26684 20130 26852 20132
rect 26684 20078 26798 20130
rect 26850 20078 26852 20130
rect 26684 20076 26852 20078
rect 26124 20020 26180 20030
rect 26124 19926 26180 19964
rect 26572 20020 26628 20030
rect 26572 19460 26628 19964
rect 26572 19394 26628 19404
rect 25340 19236 25396 19246
rect 25452 19236 25508 19246
rect 25396 19234 25508 19236
rect 25396 19182 25454 19234
rect 25506 19182 25508 19234
rect 25396 19180 25508 19182
rect 25116 19010 25172 19022
rect 25116 18958 25118 19010
rect 25170 18958 25172 19010
rect 25116 18564 25172 18958
rect 25116 18498 25172 18508
rect 24892 18274 24948 18284
rect 25340 18338 25396 19180
rect 25452 19170 25508 19180
rect 26236 19122 26292 19134
rect 26236 19070 26238 19122
rect 26290 19070 26292 19122
rect 26236 18452 26292 19070
rect 26236 18386 26292 18396
rect 26572 18564 26628 18574
rect 26572 18340 26628 18508
rect 25340 18286 25342 18338
rect 25394 18286 25396 18338
rect 24444 16046 24446 16098
rect 24498 16046 24500 16098
rect 24444 15988 24500 16046
rect 24444 15922 24500 15932
rect 24668 17556 24724 17566
rect 24668 15986 24724 17500
rect 24892 17442 24948 17454
rect 24892 17390 24894 17442
rect 24946 17390 24948 17442
rect 24892 16772 24948 17390
rect 24892 16706 24948 16716
rect 25228 16884 25284 16894
rect 25340 16884 25396 18286
rect 26460 18338 26628 18340
rect 26460 18286 26574 18338
rect 26626 18286 26628 18338
rect 26460 18284 26628 18286
rect 25788 17556 25844 17566
rect 25788 17462 25844 17500
rect 25228 16882 25396 16884
rect 25228 16830 25230 16882
rect 25282 16830 25396 16882
rect 25228 16828 25396 16830
rect 25452 17442 25508 17454
rect 25452 17390 25454 17442
rect 25506 17390 25508 17442
rect 25228 16772 25284 16828
rect 25228 16706 25284 16716
rect 25116 16100 25172 16110
rect 25452 16100 25508 17390
rect 25676 17444 25732 17454
rect 25676 17350 25732 17388
rect 26012 16772 26068 16782
rect 25788 16770 26068 16772
rect 25788 16718 26014 16770
rect 26066 16718 26068 16770
rect 25788 16716 26068 16718
rect 25676 16100 25732 16110
rect 25452 16098 25732 16100
rect 25452 16046 25678 16098
rect 25730 16046 25732 16098
rect 25452 16044 25732 16046
rect 25116 16006 25172 16044
rect 25676 16034 25732 16044
rect 25340 15988 25396 15998
rect 24668 15934 24670 15986
rect 24722 15934 24724 15986
rect 23996 15874 24164 15876
rect 23996 15822 23998 15874
rect 24050 15822 24164 15874
rect 23996 15820 24164 15822
rect 23996 15810 24052 15820
rect 24108 15316 24164 15820
rect 23548 15092 23716 15148
rect 23436 13346 23492 13356
rect 23548 12292 23604 12302
rect 23548 12198 23604 12236
rect 23212 11566 23214 11618
rect 23266 11566 23268 11618
rect 23212 11554 23268 11566
rect 23324 11282 23380 11294
rect 23324 11230 23326 11282
rect 23378 11230 23380 11282
rect 23212 11172 23268 11182
rect 22652 10498 22932 10500
rect 22652 10446 22878 10498
rect 22930 10446 22932 10498
rect 22652 10444 22932 10446
rect 20860 8530 20916 8540
rect 21756 9268 21812 9278
rect 21756 8372 21812 9212
rect 21756 8306 21812 8316
rect 19740 8260 19796 8270
rect 19628 8258 19796 8260
rect 19628 8206 19742 8258
rect 19794 8206 19796 8258
rect 19628 8204 19796 8206
rect 19740 8194 19796 8204
rect 20300 8258 20356 8270
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 17948 8034 18004 8046
rect 17948 7982 17950 8034
rect 18002 7982 18004 8034
rect 16268 7298 16324 7308
rect 16604 7362 16660 7374
rect 16604 7310 16606 7362
rect 16658 7310 16660 7362
rect 14700 6078 14702 6130
rect 14754 6078 14756 6130
rect 14700 6066 14756 6078
rect 14812 6804 14868 6814
rect 14812 6018 14868 6748
rect 16380 6804 16436 6814
rect 16380 6710 16436 6748
rect 16604 6692 16660 7310
rect 17052 7364 17108 7374
rect 17052 6692 17108 7308
rect 17948 7364 18004 7982
rect 19516 8036 19572 8046
rect 18508 7588 18564 7598
rect 18508 7494 18564 7532
rect 19180 7588 19236 7598
rect 19516 7588 19572 7980
rect 20300 8036 20356 8206
rect 20636 8260 20692 8270
rect 20636 8166 20692 8204
rect 20300 7970 20356 7980
rect 20524 8034 20580 8046
rect 20524 7982 20526 8034
rect 20578 7982 20580 8034
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19236 7532 19572 7588
rect 20412 7588 20468 7598
rect 20524 7588 20580 7982
rect 22652 8036 22708 10444
rect 22876 10434 22932 10444
rect 23100 11170 23268 11172
rect 23100 11118 23214 11170
rect 23266 11118 23268 11170
rect 23100 11116 23268 11118
rect 23100 8596 23156 11116
rect 23212 11106 23268 11116
rect 23324 10724 23380 11230
rect 23436 10724 23492 10734
rect 23324 10668 23436 10724
rect 23436 10630 23492 10668
rect 23548 10722 23604 10734
rect 23548 10670 23550 10722
rect 23602 10670 23604 10722
rect 23548 10500 23604 10670
rect 23436 10444 23604 10500
rect 23436 9380 23492 10444
rect 23548 10052 23604 10062
rect 23660 10052 23716 15092
rect 23996 14306 24052 14318
rect 23996 14254 23998 14306
rect 24050 14254 24052 14306
rect 23884 13634 23940 13646
rect 23884 13582 23886 13634
rect 23938 13582 23940 13634
rect 23884 12402 23940 13582
rect 23884 12350 23886 12402
rect 23938 12350 23940 12402
rect 23884 12338 23940 12350
rect 23996 12292 24052 14254
rect 24108 13074 24164 15260
rect 24332 14532 24388 14542
rect 24332 14438 24388 14476
rect 24668 14532 24724 15934
rect 24668 14466 24724 14476
rect 25228 15986 25396 15988
rect 25228 15934 25342 15986
rect 25394 15934 25396 15986
rect 25228 15932 25396 15934
rect 24220 14308 24276 14318
rect 24220 13636 24276 14252
rect 24668 13748 24724 13758
rect 24668 13654 24724 13692
rect 24220 13570 24276 13580
rect 24444 13636 24500 13646
rect 24108 13022 24110 13074
rect 24162 13022 24164 13074
rect 24108 13010 24164 13022
rect 24108 12292 24164 12302
rect 23996 12290 24164 12292
rect 23996 12238 24110 12290
rect 24162 12238 24164 12290
rect 23996 12236 24164 12238
rect 24108 12226 24164 12236
rect 24444 12292 24500 13580
rect 23772 12180 23828 12190
rect 23772 12086 23828 12124
rect 24332 12180 24388 12190
rect 24332 12086 24388 12124
rect 23996 12068 24052 12078
rect 23772 11956 23828 11966
rect 23772 10834 23828 11900
rect 23996 11788 24052 12012
rect 23772 10782 23774 10834
rect 23826 10782 23828 10834
rect 23772 10770 23828 10782
rect 23884 11732 24052 11788
rect 23884 10834 23940 11732
rect 24332 11172 24388 11182
rect 24444 11172 24500 12236
rect 24332 11170 24500 11172
rect 24332 11118 24334 11170
rect 24386 11118 24500 11170
rect 24332 11116 24500 11118
rect 24556 12290 24612 12302
rect 24556 12238 24558 12290
rect 24610 12238 24612 12290
rect 24332 11060 24388 11116
rect 23884 10782 23886 10834
rect 23938 10782 23940 10834
rect 23884 10770 23940 10782
rect 23996 11004 24388 11060
rect 23548 10050 23716 10052
rect 23548 9998 23550 10050
rect 23602 9998 23716 10050
rect 23548 9996 23716 9998
rect 23772 10612 23828 10622
rect 23548 9986 23604 9996
rect 23660 9828 23716 9838
rect 23772 9828 23828 10556
rect 23660 9826 23828 9828
rect 23660 9774 23662 9826
rect 23714 9774 23828 9826
rect 23660 9772 23828 9774
rect 23660 9762 23716 9772
rect 23548 9604 23604 9614
rect 23548 9602 23716 9604
rect 23548 9550 23550 9602
rect 23602 9550 23716 9602
rect 23548 9548 23716 9550
rect 23548 9538 23604 9548
rect 23436 9324 23604 9380
rect 23436 9156 23492 9166
rect 23436 9062 23492 9100
rect 22652 7970 22708 7980
rect 22764 8540 23156 8596
rect 22540 7700 22596 7710
rect 20412 7586 20580 7588
rect 20412 7534 20414 7586
rect 20466 7534 20580 7586
rect 20412 7532 20580 7534
rect 22316 7588 22372 7598
rect 18732 7476 18788 7486
rect 18732 7382 18788 7420
rect 17948 7298 18004 7308
rect 16604 6690 17108 6692
rect 16604 6638 17054 6690
rect 17106 6638 17108 6690
rect 16604 6636 17108 6638
rect 16604 6132 16660 6636
rect 17052 6626 17108 6636
rect 17724 7252 17780 7262
rect 17724 6690 17780 7196
rect 18396 7252 18452 7262
rect 18396 7158 18452 7196
rect 17724 6638 17726 6690
rect 17778 6638 17780 6690
rect 17724 6626 17780 6638
rect 19180 6692 19236 7532
rect 20412 7522 20468 7532
rect 19628 7474 19684 7486
rect 19628 7422 19630 7474
rect 19682 7422 19684 7474
rect 19292 7364 19348 7374
rect 19628 7364 19684 7422
rect 19348 7308 19684 7364
rect 19292 7270 19348 7308
rect 19180 6636 19348 6692
rect 14812 5966 14814 6018
rect 14866 5966 14868 6018
rect 14812 5954 14868 5966
rect 16044 6130 16660 6132
rect 16044 6078 16606 6130
rect 16658 6078 16660 6130
rect 16044 6076 16660 6078
rect 12348 5182 12350 5234
rect 12402 5182 12404 5234
rect 12348 5170 12404 5182
rect 15596 5236 15652 5246
rect 16044 5236 16100 6076
rect 16604 6066 16660 6076
rect 15596 5234 16100 5236
rect 15596 5182 15598 5234
rect 15650 5182 16100 5234
rect 15596 5180 16100 5182
rect 15596 5170 15652 5180
rect 8988 5124 9044 5134
rect 8764 5122 9044 5124
rect 8764 5070 8990 5122
rect 9042 5070 9044 5122
rect 8764 5068 9044 5070
rect 8988 5058 9044 5068
rect 16044 5122 16100 5180
rect 18396 5236 18452 5246
rect 16044 5070 16046 5122
rect 16098 5070 16100 5122
rect 16044 5058 16100 5070
rect 16716 5124 16772 5134
rect 16716 5030 16772 5068
rect 14364 4564 14420 4574
rect 14364 4338 14420 4508
rect 14924 4564 14980 4574
rect 14924 4470 14980 4508
rect 14364 4286 14366 4338
rect 14418 4286 14420 4338
rect 14364 4274 14420 4286
rect 12124 4116 12180 4126
rect 11676 4114 12180 4116
rect 11676 4062 12126 4114
rect 12178 4062 12180 4114
rect 11676 4060 12180 4062
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3276 3390 3278 3442
rect 3330 3390 3332 3442
rect 3276 3378 3332 3390
rect 7196 3444 7252 3454
rect 7196 800 7252 3388
rect 10108 3444 10164 3454
rect 10108 3350 10164 3388
rect 11676 800 11732 4060
rect 12124 4050 12180 4060
rect 18396 3668 18452 5180
rect 18844 5236 18900 5246
rect 18844 5142 18900 5180
rect 19180 5234 19236 5246
rect 19180 5182 19182 5234
rect 19234 5182 19236 5234
rect 19180 5124 19236 5182
rect 19180 5058 19236 5068
rect 19292 4900 19348 6636
rect 19516 5796 19572 5806
rect 19516 5346 19572 5740
rect 19516 5294 19518 5346
rect 19570 5294 19572 5346
rect 19516 5282 19572 5294
rect 19292 4806 19348 4844
rect 19628 4340 19684 7308
rect 19852 6916 19908 6926
rect 19852 6802 19908 6860
rect 22316 6916 22372 7532
rect 22540 7362 22596 7644
rect 22540 7310 22542 7362
rect 22594 7310 22596 7362
rect 22540 7298 22596 7310
rect 19852 6750 19854 6802
rect 19906 6750 19908 6802
rect 19852 6738 19908 6750
rect 22204 6804 22260 6814
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 22204 5906 22260 6748
rect 22316 6130 22372 6860
rect 22316 6078 22318 6130
rect 22370 6078 22372 6130
rect 22316 6066 22372 6078
rect 22540 6020 22596 6030
rect 22764 6020 22820 8540
rect 22988 8370 23044 8382
rect 23548 8372 23604 9324
rect 22988 8318 22990 8370
rect 23042 8318 23044 8370
rect 22988 8260 23044 8318
rect 22988 8194 23044 8204
rect 23436 8316 23604 8372
rect 23212 8148 23268 8158
rect 22988 8034 23044 8046
rect 22988 7982 22990 8034
rect 23042 7982 23044 8034
rect 22988 7474 23044 7982
rect 23100 8036 23156 8046
rect 23100 7942 23156 7980
rect 23100 7700 23156 7710
rect 23212 7700 23268 8092
rect 23156 7644 23268 7700
rect 23324 8034 23380 8046
rect 23324 7982 23326 8034
rect 23378 7982 23380 8034
rect 23324 7812 23380 7982
rect 23324 7698 23380 7756
rect 23324 7646 23326 7698
rect 23378 7646 23380 7698
rect 23100 7606 23156 7644
rect 23324 7634 23380 7646
rect 23436 7588 23492 8316
rect 23548 8148 23604 8158
rect 23548 8054 23604 8092
rect 23548 7588 23604 7598
rect 23492 7586 23604 7588
rect 23492 7534 23550 7586
rect 23602 7534 23604 7586
rect 23492 7532 23604 7534
rect 23436 7494 23492 7532
rect 23548 7522 23604 7532
rect 22988 7422 22990 7474
rect 23042 7422 23044 7474
rect 22988 6804 23044 7422
rect 23212 7476 23268 7486
rect 23212 7382 23268 7420
rect 22988 6738 23044 6748
rect 22988 6132 23044 6142
rect 22540 5926 22596 5964
rect 22652 6018 22820 6020
rect 22652 5966 22766 6018
rect 22818 5966 22820 6018
rect 22652 5964 22820 5966
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 21308 5236 21364 5246
rect 20748 5234 21364 5236
rect 20748 5182 21310 5234
rect 21362 5182 21364 5234
rect 20748 5180 21364 5182
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20748 4450 20804 5180
rect 21308 5170 21364 5180
rect 21644 5124 21700 5134
rect 22204 5124 22260 5854
rect 22428 5796 22484 5806
rect 22428 5702 22484 5740
rect 22428 5234 22484 5246
rect 22428 5182 22430 5234
rect 22482 5182 22484 5234
rect 22316 5124 22372 5134
rect 22204 5122 22372 5124
rect 22204 5070 22318 5122
rect 22370 5070 22372 5122
rect 22204 5068 22372 5070
rect 21644 5030 21700 5068
rect 22316 5058 22372 5068
rect 22428 5124 22484 5182
rect 22652 5236 22708 5964
rect 22764 5954 22820 5964
rect 22876 6020 22932 6030
rect 22428 5058 22484 5068
rect 22540 5124 22596 5134
rect 22652 5124 22708 5180
rect 22540 5122 22708 5124
rect 22540 5070 22542 5122
rect 22594 5070 22708 5122
rect 22540 5068 22708 5070
rect 22764 5124 22820 5134
rect 22876 5124 22932 5964
rect 22764 5122 22932 5124
rect 22764 5070 22766 5122
rect 22818 5070 22932 5122
rect 22764 5068 22932 5070
rect 22988 5122 23044 6076
rect 23660 6132 23716 9548
rect 23772 9156 23828 9166
rect 23996 9156 24052 11004
rect 23772 9154 24052 9156
rect 23772 9102 23774 9154
rect 23826 9102 24052 9154
rect 23772 9100 24052 9102
rect 24108 10722 24164 10734
rect 24108 10670 24110 10722
rect 24162 10670 24164 10722
rect 23772 7588 23828 9100
rect 23772 7522 23828 7532
rect 24108 7476 24164 10670
rect 24220 10724 24276 10734
rect 24220 10630 24276 10668
rect 24556 8148 24612 12238
rect 24668 12180 24724 12190
rect 24668 12086 24724 12124
rect 25228 11956 25284 15932
rect 25340 15922 25396 15932
rect 25564 15876 25620 15886
rect 25788 15876 25844 16716
rect 26012 16706 26068 16716
rect 25564 15874 25844 15876
rect 25564 15822 25566 15874
rect 25618 15822 25844 15874
rect 25564 15820 25844 15822
rect 25564 15810 25620 15820
rect 25340 15764 25396 15774
rect 25340 14308 25396 15708
rect 26012 14532 26068 14542
rect 26012 14438 26068 14476
rect 25340 14242 25396 14252
rect 26124 14308 26180 14318
rect 26124 14214 26180 14252
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 25788 13746 25844 13758
rect 25788 13694 25790 13746
rect 25842 13694 25844 13746
rect 25340 13636 25396 13646
rect 25340 13542 25396 13580
rect 25788 13636 25844 13694
rect 25788 13570 25844 13580
rect 26012 13746 26068 13758
rect 26012 13694 26014 13746
rect 26066 13694 26068 13746
rect 26012 13300 26068 13694
rect 26348 13746 26404 14254
rect 26348 13694 26350 13746
rect 26402 13694 26404 13746
rect 26348 13682 26404 13694
rect 26124 13636 26180 13646
rect 26124 13542 26180 13580
rect 26012 13244 26404 13300
rect 26124 12962 26180 12974
rect 26124 12910 26126 12962
rect 26178 12910 26180 12962
rect 26124 12852 26180 12910
rect 26348 12962 26404 13244
rect 26348 12910 26350 12962
rect 26402 12910 26404 12962
rect 26348 12898 26404 12910
rect 25228 11890 25284 11900
rect 25788 12796 26124 12852
rect 25788 12178 25844 12796
rect 26124 12786 26180 12796
rect 25788 12126 25790 12178
rect 25842 12126 25844 12178
rect 25788 11844 25844 12126
rect 25788 11778 25844 11788
rect 25900 12180 25956 12190
rect 25900 11844 25956 12124
rect 26124 11844 26180 11854
rect 25900 11788 26124 11844
rect 25900 11282 25956 11788
rect 26124 11778 26180 11788
rect 25900 11230 25902 11282
rect 25954 11230 25956 11282
rect 25900 11218 25956 11230
rect 26348 11284 26404 11294
rect 26236 11170 26292 11182
rect 26236 11118 26238 11170
rect 26290 11118 26292 11170
rect 25228 10724 25284 10734
rect 25228 10630 25284 10668
rect 25564 10610 25620 10622
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 25564 10500 25620 10558
rect 26012 10500 26068 10510
rect 25564 10498 26068 10500
rect 25564 10446 26014 10498
rect 26066 10446 26068 10498
rect 25564 10444 26068 10446
rect 26012 10164 26068 10444
rect 26236 10276 26292 11118
rect 26236 10210 26292 10220
rect 26012 10098 26068 10108
rect 26236 9268 26292 9278
rect 26348 9268 26404 11228
rect 26460 11172 26516 18284
rect 26572 18274 26628 18284
rect 26796 14980 26852 20076
rect 27132 18564 27188 18574
rect 27132 18470 27188 18508
rect 26908 18450 26964 18462
rect 26908 18398 26910 18450
rect 26962 18398 26964 18450
rect 26908 15148 26964 18398
rect 27020 18452 27076 18462
rect 27020 18358 27076 18396
rect 27468 15148 27524 21980
rect 27804 21924 27860 22316
rect 28028 22306 28084 22316
rect 27580 21868 27860 21924
rect 27580 21810 27636 21868
rect 27580 21758 27582 21810
rect 27634 21758 27636 21810
rect 27580 21746 27636 21758
rect 27580 19012 27636 19022
rect 27580 18450 27636 18956
rect 27580 18398 27582 18450
rect 27634 18398 27636 18450
rect 27580 18386 27636 18398
rect 28252 17444 28308 26852
rect 28588 26180 28644 28476
rect 30044 28532 30100 36204
rect 30156 36194 30212 36204
rect 30604 35810 30660 35822
rect 30604 35758 30606 35810
rect 30658 35758 30660 35810
rect 30156 35698 30212 35710
rect 30156 35646 30158 35698
rect 30210 35646 30212 35698
rect 30156 35588 30212 35646
rect 30156 35364 30212 35532
rect 30156 35308 30436 35364
rect 30156 35028 30212 35038
rect 30156 34934 30212 34972
rect 30044 28466 30100 28476
rect 30268 30100 30324 30110
rect 30268 29986 30324 30044
rect 30268 29934 30270 29986
rect 30322 29934 30324 29986
rect 29708 28196 29764 28206
rect 29036 26964 29092 26974
rect 28588 26114 28644 26124
rect 28924 26628 28980 26638
rect 28476 25284 28532 25294
rect 28532 25228 28644 25284
rect 28476 25190 28532 25228
rect 28588 25172 28644 25228
rect 28588 25116 28756 25172
rect 28588 24948 28644 24958
rect 28364 24836 28420 24846
rect 28364 24742 28420 24780
rect 28588 24834 28644 24892
rect 28588 24782 28590 24834
rect 28642 24782 28644 24834
rect 28588 24770 28644 24782
rect 28700 24276 28756 25116
rect 28924 24836 28980 26572
rect 29036 26402 29092 26908
rect 29036 26350 29038 26402
rect 29090 26350 29092 26402
rect 29036 26338 29092 26350
rect 29148 26852 29204 26862
rect 29148 25394 29204 26796
rect 29708 25620 29764 28140
rect 30268 26404 30324 29934
rect 30380 28420 30436 35308
rect 30604 34916 30660 35758
rect 30604 34850 30660 34860
rect 30604 34692 30660 34702
rect 30604 34598 30660 34636
rect 30604 34020 30660 34030
rect 30604 33926 30660 33964
rect 30828 32340 30884 37324
rect 31836 36372 31892 36382
rect 31724 36316 31836 36372
rect 30940 35698 30996 35710
rect 30940 35646 30942 35698
rect 30994 35646 30996 35698
rect 30940 34804 30996 35646
rect 31612 35700 31668 35710
rect 31612 35606 31668 35644
rect 31052 35028 31108 35038
rect 31052 34914 31108 34972
rect 31724 35026 31780 36316
rect 31836 36306 31892 36316
rect 32172 35698 32228 38612
rect 32620 35924 32676 35934
rect 32620 35830 32676 35868
rect 32396 35810 32452 35822
rect 32396 35758 32398 35810
rect 32450 35758 32452 35810
rect 32172 35646 32174 35698
rect 32226 35646 32228 35698
rect 32172 35634 32228 35646
rect 32284 35700 32340 35710
rect 31724 34974 31726 35026
rect 31778 34974 31780 35026
rect 31724 34962 31780 34974
rect 31052 34862 31054 34914
rect 31106 34862 31108 34914
rect 31052 34850 31108 34862
rect 31276 34916 31332 34926
rect 30940 34738 30996 34748
rect 31276 34802 31332 34860
rect 31276 34750 31278 34802
rect 31330 34750 31332 34802
rect 31276 34738 31332 34750
rect 31948 34914 32004 34926
rect 31948 34862 31950 34914
rect 32002 34862 32004 34914
rect 31948 34804 32004 34862
rect 31948 34738 32004 34748
rect 31612 33348 31668 33358
rect 30828 32274 30884 32284
rect 31052 33346 31668 33348
rect 31052 33294 31614 33346
rect 31666 33294 31668 33346
rect 31052 33292 31668 33294
rect 31052 31890 31108 33292
rect 31612 33282 31668 33292
rect 31052 31838 31054 31890
rect 31106 31838 31108 31890
rect 31052 31826 31108 31838
rect 31164 33124 31220 33134
rect 31164 32004 31220 33068
rect 32284 32788 32340 35644
rect 32396 34916 32452 35758
rect 32396 34850 32452 34860
rect 32620 34914 32676 34926
rect 32620 34862 32622 34914
rect 32674 34862 32676 34914
rect 32620 34692 32676 34862
rect 32956 34914 33012 38612
rect 33180 38164 33236 39006
rect 33516 38164 33572 38174
rect 33068 38108 33516 38164
rect 33068 38050 33124 38108
rect 33516 38098 33572 38108
rect 33068 37998 33070 38050
rect 33122 37998 33124 38050
rect 33068 37986 33124 37998
rect 33740 37940 33796 37950
rect 33740 37938 33908 37940
rect 33740 37886 33742 37938
rect 33794 37886 33908 37938
rect 33740 37884 33908 37886
rect 33740 37874 33796 37884
rect 33180 35700 33236 35710
rect 33180 35606 33236 35644
rect 33516 35140 33572 35150
rect 32956 34862 32958 34914
rect 33010 34862 33012 34914
rect 32956 34850 33012 34862
rect 33404 34916 33460 34926
rect 33404 34802 33460 34860
rect 33404 34750 33406 34802
rect 33458 34750 33460 34802
rect 33404 34738 33460 34750
rect 32620 34626 32676 34636
rect 33404 34356 33460 34366
rect 33516 34356 33572 35084
rect 33852 35138 33908 37884
rect 34076 35810 34132 35822
rect 34076 35758 34078 35810
rect 34130 35758 34132 35810
rect 33852 35086 33854 35138
rect 33906 35086 33908 35138
rect 33852 35074 33908 35086
rect 33964 35698 34020 35710
rect 33964 35646 33966 35698
rect 34018 35646 34020 35698
rect 33404 34354 33572 34356
rect 33404 34302 33406 34354
rect 33458 34302 33572 34354
rect 33404 34300 33572 34302
rect 33404 34290 33460 34300
rect 33292 34244 33348 34254
rect 32396 34020 32452 34030
rect 32396 33460 32452 33964
rect 32396 33346 32452 33404
rect 32844 33460 32900 33470
rect 32844 33366 32900 33404
rect 32396 33294 32398 33346
rect 32450 33294 32452 33346
rect 32396 33282 32452 33294
rect 32284 32732 32452 32788
rect 31724 32004 31780 32014
rect 30828 31554 30884 31566
rect 30828 31502 30830 31554
rect 30882 31502 30884 31554
rect 30492 31444 30548 31454
rect 30492 31218 30548 31388
rect 30828 31220 30884 31502
rect 30492 31166 30494 31218
rect 30546 31166 30548 31218
rect 30492 29540 30548 31166
rect 30604 31164 30884 31220
rect 31052 31554 31108 31566
rect 31052 31502 31054 31554
rect 31106 31502 31108 31554
rect 31052 31218 31108 31502
rect 31052 31166 31054 31218
rect 31106 31166 31108 31218
rect 30604 29764 30660 31164
rect 31052 31154 31108 31166
rect 30828 30994 30884 31006
rect 30828 30942 30830 30994
rect 30882 30942 30884 30994
rect 30828 30884 30884 30942
rect 30828 29764 30884 30828
rect 31164 29764 31220 31948
rect 31388 32002 31780 32004
rect 31388 31950 31726 32002
rect 31778 31950 31780 32002
rect 31388 31948 31780 31950
rect 31388 31778 31444 31948
rect 31724 31938 31780 31948
rect 31388 31726 31390 31778
rect 31442 31726 31444 31778
rect 31388 31714 31444 31726
rect 31724 31780 31780 31790
rect 31612 31666 31668 31678
rect 31612 31614 31614 31666
rect 31666 31614 31668 31666
rect 31612 31444 31668 31614
rect 31724 31666 31780 31724
rect 32284 31780 32340 31790
rect 32284 31686 32340 31724
rect 31724 31614 31726 31666
rect 31778 31614 31780 31666
rect 31724 31602 31780 31614
rect 31612 31378 31668 31388
rect 31276 31220 31332 31230
rect 31276 31218 31556 31220
rect 31276 31166 31278 31218
rect 31330 31166 31556 31218
rect 31276 31164 31556 31166
rect 31276 30996 31332 31164
rect 31500 31108 31556 31164
rect 31836 31108 31892 31118
rect 31500 31106 31892 31108
rect 31500 31054 31838 31106
rect 31890 31054 31892 31106
rect 31500 31052 31892 31054
rect 31276 30930 31332 30940
rect 31388 30996 31444 31006
rect 31388 30994 31668 30996
rect 31388 30942 31390 30994
rect 31442 30942 31668 30994
rect 31388 30940 31668 30942
rect 31388 30930 31444 30940
rect 31276 30436 31332 30446
rect 31276 30434 31556 30436
rect 31276 30382 31278 30434
rect 31330 30382 31556 30434
rect 31276 30380 31556 30382
rect 31276 30370 31332 30380
rect 31388 30212 31444 30222
rect 31388 30118 31444 30156
rect 31276 29988 31332 29998
rect 31276 29894 31332 29932
rect 30828 29708 30996 29764
rect 31164 29708 31444 29764
rect 30604 29698 30660 29708
rect 30716 29540 30772 29550
rect 30492 29538 30772 29540
rect 30492 29486 30718 29538
rect 30770 29486 30772 29538
rect 30492 29484 30772 29486
rect 30492 28420 30548 28430
rect 30380 28364 30492 28420
rect 30492 28326 30548 28364
rect 30604 28196 30660 29484
rect 30716 29474 30772 29484
rect 30828 29538 30884 29550
rect 30828 29486 30830 29538
rect 30882 29486 30884 29538
rect 30828 29428 30884 29486
rect 30828 29362 30884 29372
rect 30940 29316 30996 29708
rect 31052 29652 31108 29662
rect 31052 29650 31332 29652
rect 31052 29598 31054 29650
rect 31106 29598 31332 29650
rect 31052 29596 31332 29598
rect 31052 29586 31108 29596
rect 31276 29538 31332 29596
rect 31276 29486 31278 29538
rect 31330 29486 31332 29538
rect 31276 29474 31332 29486
rect 31388 29316 31444 29708
rect 31500 29650 31556 30380
rect 31612 30212 31668 30940
rect 31612 30146 31668 30156
rect 31836 29988 31892 31052
rect 31500 29598 31502 29650
rect 31554 29598 31556 29650
rect 31500 29586 31556 29598
rect 31612 29932 31892 29988
rect 31948 29988 32004 29998
rect 30940 29260 31108 29316
rect 30940 28530 30996 28542
rect 30940 28478 30942 28530
rect 30994 28478 30996 28530
rect 30492 28140 30660 28196
rect 30716 28418 30772 28430
rect 30716 28366 30718 28418
rect 30770 28366 30772 28418
rect 30268 26338 30324 26348
rect 30380 27972 30436 27982
rect 29820 26290 29876 26302
rect 29820 26238 29822 26290
rect 29874 26238 29876 26290
rect 29820 26180 29876 26238
rect 29820 26114 29876 26124
rect 30268 26180 30324 26190
rect 30268 26086 30324 26124
rect 29708 25564 30100 25620
rect 29372 25508 29428 25518
rect 29372 25414 29428 25452
rect 29148 25342 29150 25394
rect 29202 25342 29204 25394
rect 29148 25330 29204 25342
rect 29932 25396 29988 25406
rect 29932 25302 29988 25340
rect 29596 25004 29988 25060
rect 29148 24948 29204 24958
rect 29596 24948 29652 25004
rect 29148 24946 29652 24948
rect 29148 24894 29150 24946
rect 29202 24894 29652 24946
rect 29148 24892 29652 24894
rect 29148 24882 29204 24892
rect 28924 24770 28980 24780
rect 29708 24836 29764 24846
rect 29708 24742 29764 24780
rect 29036 24724 29092 24734
rect 29596 24724 29652 24734
rect 29036 24630 29092 24668
rect 29372 24722 29652 24724
rect 29372 24670 29598 24722
rect 29650 24670 29652 24722
rect 29372 24668 29652 24670
rect 28924 24500 28980 24510
rect 29372 24500 29428 24668
rect 29596 24658 29652 24668
rect 28924 24498 29428 24500
rect 28924 24446 28926 24498
rect 28978 24446 29428 24498
rect 28924 24444 29428 24446
rect 29484 24498 29540 24510
rect 29484 24446 29486 24498
rect 29538 24446 29540 24498
rect 28924 24434 28980 24444
rect 29484 24388 29540 24446
rect 29036 24332 29540 24388
rect 29036 24276 29092 24332
rect 28700 24220 29092 24276
rect 29932 24050 29988 25004
rect 29932 23998 29934 24050
rect 29986 23998 29988 24050
rect 29932 23986 29988 23998
rect 29260 23938 29316 23950
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 28588 23716 28644 23726
rect 29260 23716 29316 23886
rect 28588 23714 29316 23716
rect 28588 23662 28590 23714
rect 28642 23662 29316 23714
rect 28588 23660 29316 23662
rect 28588 23044 28644 23660
rect 28588 22978 28644 22988
rect 29260 22708 29316 23660
rect 29260 22642 29316 22652
rect 29148 22484 29204 22494
rect 29148 20916 29204 22428
rect 29932 22484 29988 22494
rect 30044 22484 30100 25564
rect 30380 25508 30436 27916
rect 30492 27074 30548 28140
rect 30716 27636 30772 28366
rect 30828 28420 30884 28430
rect 30940 28420 30996 28478
rect 30884 28364 30996 28420
rect 31052 28530 31108 29260
rect 31052 28478 31054 28530
rect 31106 28478 31108 28530
rect 30828 28354 30884 28364
rect 30716 27580 30884 27636
rect 30492 27022 30494 27074
rect 30546 27022 30548 27074
rect 30492 26740 30548 27022
rect 30716 27188 30772 27198
rect 30604 26964 30660 27002
rect 30604 26898 30660 26908
rect 30716 26962 30772 27132
rect 30716 26910 30718 26962
rect 30770 26910 30772 26962
rect 30716 26898 30772 26910
rect 30828 26962 30884 27580
rect 31052 27300 31108 28478
rect 31276 29260 31444 29316
rect 31276 27972 31332 29260
rect 31388 28756 31444 28766
rect 31388 28642 31444 28700
rect 31388 28590 31390 28642
rect 31442 28590 31444 28642
rect 31388 28578 31444 28590
rect 31276 27878 31332 27916
rect 31612 27748 31668 29932
rect 31948 29894 32004 29932
rect 31724 29764 31780 29774
rect 31724 29650 31780 29708
rect 31724 29598 31726 29650
rect 31778 29598 31780 29650
rect 31724 29586 31780 29598
rect 32172 29428 32228 29438
rect 32172 29334 32228 29372
rect 31836 29204 31892 29214
rect 31836 29202 32116 29204
rect 31836 29150 31838 29202
rect 31890 29150 32116 29202
rect 31836 29148 32116 29150
rect 31836 29138 31892 29148
rect 32060 28756 32116 29148
rect 32172 28756 32228 28766
rect 32060 28754 32228 28756
rect 32060 28702 32174 28754
rect 32226 28702 32228 28754
rect 32060 28700 32228 28702
rect 32172 28690 32228 28700
rect 31052 27234 31108 27244
rect 31164 27692 31668 27748
rect 31724 28532 31780 28542
rect 30828 26910 30830 26962
rect 30882 26910 30884 26962
rect 30828 26898 30884 26910
rect 31164 26908 31220 27692
rect 31276 27076 31332 27086
rect 31276 27074 31668 27076
rect 31276 27022 31278 27074
rect 31330 27022 31668 27074
rect 31276 27020 31668 27022
rect 31276 27010 31332 27020
rect 31052 26852 31220 26908
rect 31612 26964 31668 27020
rect 31500 26852 31556 26862
rect 30492 26684 30996 26740
rect 30940 26514 30996 26684
rect 30940 26462 30942 26514
rect 30994 26462 30996 26514
rect 30940 26450 30996 26462
rect 30828 26292 30884 26302
rect 30156 25452 30436 25508
rect 30492 25508 30548 25518
rect 30156 24724 30212 25452
rect 30492 25396 30548 25452
rect 30380 25340 30548 25396
rect 30380 25282 30436 25340
rect 30380 25230 30382 25282
rect 30434 25230 30436 25282
rect 30380 25218 30436 25230
rect 30268 24948 30324 24958
rect 30268 24854 30324 24892
rect 30604 24836 30660 24846
rect 30604 24724 30660 24780
rect 30716 24724 30772 24734
rect 30156 24668 30324 24724
rect 30604 24722 30772 24724
rect 30604 24670 30718 24722
rect 30770 24670 30772 24722
rect 30604 24668 30772 24670
rect 29932 22482 30100 22484
rect 29932 22430 29934 22482
rect 29986 22430 30100 22482
rect 29932 22428 30100 22430
rect 29932 22418 29988 22428
rect 29484 22370 29540 22382
rect 29484 22318 29486 22370
rect 29538 22318 29540 22370
rect 29484 22148 29540 22318
rect 29484 22082 29540 22092
rect 30044 21700 30100 22428
rect 29932 20916 29988 20926
rect 29148 20860 29428 20916
rect 29148 20692 29204 20702
rect 29148 20598 29204 20636
rect 29260 20578 29316 20590
rect 29260 20526 29262 20578
rect 29314 20526 29316 20578
rect 29260 19236 29316 20526
rect 29148 19180 29316 19236
rect 29372 19236 29428 20860
rect 29932 20822 29988 20860
rect 30044 20692 30100 21644
rect 30268 20692 30324 24668
rect 30716 24658 30772 24668
rect 30380 22148 30436 22158
rect 30380 21476 30436 22092
rect 30828 22148 30884 26236
rect 31052 25172 31108 26852
rect 31388 26850 31556 26852
rect 31388 26798 31502 26850
rect 31554 26798 31556 26850
rect 31388 26796 31556 26798
rect 31164 26402 31220 26414
rect 31164 26350 31166 26402
rect 31218 26350 31220 26402
rect 31164 25732 31220 26350
rect 31388 26290 31444 26796
rect 31500 26786 31556 26796
rect 31388 26238 31390 26290
rect 31442 26238 31444 26290
rect 31388 26226 31444 26238
rect 31612 26290 31668 26908
rect 31724 26962 31780 28476
rect 31836 27300 31892 27310
rect 31836 27074 31892 27244
rect 32284 27188 32340 27198
rect 32284 27094 32340 27132
rect 31836 27022 31838 27074
rect 31890 27022 31892 27074
rect 31836 27010 31892 27022
rect 31948 27076 32004 27086
rect 31724 26910 31726 26962
rect 31778 26910 31780 26962
rect 31724 26898 31780 26910
rect 31948 26908 32004 27020
rect 31612 26238 31614 26290
rect 31666 26238 31668 26290
rect 31612 26226 31668 26238
rect 31836 26852 32004 26908
rect 31164 25666 31220 25676
rect 31276 26180 31332 26190
rect 31276 25506 31332 26124
rect 31724 26178 31780 26190
rect 31724 26126 31726 26178
rect 31778 26126 31780 26178
rect 31724 25620 31780 26126
rect 31724 25554 31780 25564
rect 31276 25454 31278 25506
rect 31330 25454 31332 25506
rect 31276 25284 31332 25454
rect 31276 25218 31332 25228
rect 31052 25116 31220 25172
rect 31164 25060 31220 25116
rect 31164 25004 31332 25060
rect 31052 24948 31108 24958
rect 30828 22082 30884 22092
rect 30940 24892 31052 24948
rect 30380 21410 30436 21420
rect 30716 21476 30772 21486
rect 30940 21476 30996 24892
rect 31052 24882 31108 24892
rect 30716 21474 30996 21476
rect 30716 21422 30718 21474
rect 30770 21422 30996 21474
rect 30716 21420 30996 21422
rect 31164 22484 31220 22494
rect 30044 20626 30100 20636
rect 30156 20636 30324 20692
rect 30380 20804 30436 20814
rect 30716 20804 30772 21420
rect 30380 20802 30772 20804
rect 30380 20750 30382 20802
rect 30434 20750 30772 20802
rect 30380 20748 30772 20750
rect 31164 20802 31220 22428
rect 31164 20750 31166 20802
rect 31218 20750 31220 20802
rect 29484 20578 29540 20590
rect 29484 20526 29486 20578
rect 29538 20526 29540 20578
rect 29484 19908 29540 20526
rect 29484 19842 29540 19852
rect 30156 19796 30212 20636
rect 30380 20356 30436 20748
rect 31164 20738 31220 20750
rect 30828 20692 30884 20702
rect 30828 20598 30884 20636
rect 30940 20580 30996 20590
rect 30940 20578 31108 20580
rect 30940 20526 30942 20578
rect 30994 20526 31108 20578
rect 30940 20524 31108 20526
rect 30940 20514 30996 20524
rect 30268 20300 30436 20356
rect 30268 20020 30324 20300
rect 30268 19926 30324 19964
rect 30492 20130 30548 20142
rect 30492 20078 30494 20130
rect 30546 20078 30548 20130
rect 30492 19796 30548 20078
rect 30156 19740 30436 19796
rect 28476 19124 28532 19134
rect 28476 19010 28532 19068
rect 28476 18958 28478 19010
rect 28530 18958 28532 19010
rect 28476 18946 28532 18958
rect 29036 19012 29092 19022
rect 29036 18918 29092 18956
rect 29148 17892 29204 19180
rect 29260 19012 29316 19022
rect 29260 18918 29316 18956
rect 29148 17836 29316 17892
rect 29148 17666 29204 17678
rect 29148 17614 29150 17666
rect 29202 17614 29204 17666
rect 28140 16772 28196 16782
rect 28252 16772 28308 17388
rect 28140 16770 28308 16772
rect 28140 16718 28142 16770
rect 28194 16718 28308 16770
rect 28140 16716 28308 16718
rect 28588 17444 28644 17454
rect 29148 17444 29204 17614
rect 28588 17442 29204 17444
rect 28588 17390 28590 17442
rect 28642 17390 29204 17442
rect 28588 17388 29204 17390
rect 28140 16706 28196 16716
rect 28476 15316 28532 15326
rect 28588 15316 28644 17388
rect 28812 15988 28868 15998
rect 28812 15538 28868 15932
rect 29260 15764 29316 17836
rect 29260 15698 29316 15708
rect 29372 15540 29428 19180
rect 30268 19236 30324 19246
rect 30268 19142 30324 19180
rect 29820 19012 29876 19022
rect 29820 18918 29876 18956
rect 30380 18788 30436 19740
rect 30492 19730 30548 19740
rect 30828 20020 30884 20030
rect 30828 19908 30884 19964
rect 30940 19908 30996 19918
rect 30828 19906 30996 19908
rect 30828 19854 30942 19906
rect 30994 19854 30996 19906
rect 30828 19852 30996 19854
rect 30268 18732 30436 18788
rect 29932 18340 29988 18350
rect 29932 17778 29988 18284
rect 29932 17726 29934 17778
rect 29986 17726 29988 17778
rect 29932 17714 29988 17726
rect 28812 15486 28814 15538
rect 28866 15486 28868 15538
rect 28812 15474 28868 15486
rect 29036 15484 29428 15540
rect 30268 17108 30324 18732
rect 28532 15260 28644 15316
rect 28476 15222 28532 15260
rect 26908 15092 27076 15148
rect 26796 14914 26852 14924
rect 26572 13748 26628 13758
rect 26628 13692 26964 13748
rect 26572 13654 26628 13692
rect 26684 13300 26740 13310
rect 26684 12962 26740 13244
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26572 12740 26628 12750
rect 26572 12646 26628 12684
rect 26684 11844 26740 12910
rect 26572 11396 26628 11406
rect 26684 11396 26740 11788
rect 26572 11394 26740 11396
rect 26572 11342 26574 11394
rect 26626 11342 26740 11394
rect 26572 11340 26740 11342
rect 26908 12068 26964 13692
rect 27020 13300 27076 15092
rect 27020 13234 27076 13244
rect 27244 15092 27524 15148
rect 27132 12852 27188 12862
rect 27132 12738 27188 12796
rect 27132 12686 27134 12738
rect 27186 12686 27188 12738
rect 27132 12404 27188 12686
rect 27132 12338 27188 12348
rect 26572 11330 26628 11340
rect 26796 11284 26852 11294
rect 26796 11190 26852 11228
rect 26460 11116 26628 11172
rect 26572 10948 26628 11116
rect 26572 10892 26852 10948
rect 26236 9266 26740 9268
rect 26236 9214 26238 9266
rect 26290 9214 26740 9266
rect 26236 9212 26740 9214
rect 26236 9202 26292 9212
rect 26124 8930 26180 8942
rect 26124 8878 26126 8930
rect 26178 8878 26180 8930
rect 26124 8820 26180 8878
rect 25228 8764 26628 8820
rect 25228 8258 25284 8764
rect 25340 8596 25396 8606
rect 25340 8370 25396 8540
rect 25340 8318 25342 8370
rect 25394 8318 25396 8370
rect 25340 8306 25396 8318
rect 26236 8372 26292 8382
rect 26236 8278 26292 8316
rect 25228 8206 25230 8258
rect 25282 8206 25284 8258
rect 25228 8194 25284 8206
rect 25452 8258 25508 8270
rect 25452 8206 25454 8258
rect 25506 8206 25508 8258
rect 24556 8082 24612 8092
rect 24780 8146 24836 8158
rect 24780 8094 24782 8146
rect 24834 8094 24836 8146
rect 24780 8036 24836 8094
rect 25452 8148 25508 8206
rect 26012 8258 26068 8270
rect 26012 8206 26014 8258
rect 26066 8206 26068 8258
rect 25452 8082 25508 8092
rect 25788 8146 25844 8158
rect 25788 8094 25790 8146
rect 25842 8094 25844 8146
rect 24780 7970 24836 7980
rect 25004 8034 25060 8046
rect 25004 7982 25006 8034
rect 25058 7982 25060 8034
rect 25004 7812 25060 7982
rect 25004 7746 25060 7756
rect 24108 7420 24612 7476
rect 23884 6804 23940 6814
rect 23884 6578 23940 6748
rect 23884 6526 23886 6578
rect 23938 6526 23940 6578
rect 23884 6514 23940 6526
rect 24220 6468 24276 6478
rect 23660 6066 23716 6076
rect 24108 6412 24220 6468
rect 24108 6130 24164 6412
rect 24220 6374 24276 6412
rect 24108 6078 24110 6130
rect 24162 6078 24164 6130
rect 24108 6066 24164 6078
rect 24220 6132 24276 6142
rect 24220 6038 24276 6076
rect 24444 6132 24500 6142
rect 24444 6038 24500 6076
rect 24556 5908 24612 7420
rect 25452 7364 25508 7374
rect 25788 7364 25844 8094
rect 26012 8148 26068 8206
rect 26012 8082 26068 8092
rect 26460 8146 26516 8158
rect 26460 8094 26462 8146
rect 26514 8094 26516 8146
rect 26348 8036 26404 8046
rect 26348 7942 26404 7980
rect 25900 7812 25956 7822
rect 26460 7812 26516 8094
rect 25956 7756 26516 7812
rect 25900 7698 25956 7756
rect 25900 7646 25902 7698
rect 25954 7646 25956 7698
rect 25900 7634 25956 7646
rect 26236 7476 26292 7486
rect 26236 7382 26292 7420
rect 25452 7362 25844 7364
rect 25452 7310 25454 7362
rect 25506 7310 25844 7362
rect 25452 7308 25844 7310
rect 26572 7362 26628 8764
rect 26684 8258 26740 9212
rect 26684 8206 26686 8258
rect 26738 8206 26740 8258
rect 26684 8194 26740 8206
rect 26572 7310 26574 7362
rect 26626 7310 26628 7362
rect 25452 7028 25508 7308
rect 26572 7298 26628 7310
rect 25452 6962 25508 6972
rect 26796 6692 26852 10892
rect 26908 10612 26964 12012
rect 27244 11732 27300 15092
rect 27580 14980 27636 14990
rect 27356 13636 27412 13646
rect 27356 13542 27412 13580
rect 27132 11676 27300 11732
rect 27132 11508 27188 11676
rect 27580 11508 27636 14924
rect 28252 12404 28308 12414
rect 28252 12310 28308 12348
rect 27916 11508 27972 11518
rect 27132 11452 27300 11508
rect 27020 11396 27076 11406
rect 27020 11302 27076 11340
rect 26908 10610 27076 10612
rect 26908 10558 26910 10610
rect 26962 10558 27076 10610
rect 26908 10556 27076 10558
rect 26908 10546 26964 10556
rect 27020 7364 27076 10556
rect 27132 10276 27188 10286
rect 27132 9828 27188 10220
rect 27244 10050 27300 11452
rect 27580 11506 27972 11508
rect 27580 11454 27918 11506
rect 27970 11454 27972 11506
rect 27580 11452 27972 11454
rect 27356 11396 27412 11406
rect 27580 11396 27636 11452
rect 27916 11442 27972 11452
rect 27356 11394 27636 11396
rect 27356 11342 27358 11394
rect 27410 11342 27636 11394
rect 27356 11340 27636 11342
rect 27356 11330 27412 11340
rect 27356 11172 27412 11182
rect 27356 11170 27636 11172
rect 27356 11118 27358 11170
rect 27410 11118 27636 11170
rect 27356 11116 27636 11118
rect 27356 11106 27412 11116
rect 27580 10722 27636 11116
rect 27580 10670 27582 10722
rect 27634 10670 27636 10722
rect 27580 10658 27636 10670
rect 27244 9998 27246 10050
rect 27298 9998 27300 10050
rect 27244 9986 27300 9998
rect 27132 9734 27188 9772
rect 27244 9604 27300 9614
rect 27244 9602 27412 9604
rect 27244 9550 27246 9602
rect 27298 9550 27412 9602
rect 27244 9548 27412 9550
rect 27244 9538 27300 9548
rect 27244 8372 27300 8382
rect 27244 8278 27300 8316
rect 27020 7298 27076 7308
rect 27020 7028 27076 7038
rect 26796 6636 26964 6692
rect 26684 6466 26740 6478
rect 26684 6414 26686 6466
rect 26738 6414 26740 6466
rect 26684 6132 26740 6414
rect 26684 6066 26740 6076
rect 24556 5814 24612 5852
rect 24332 5794 24388 5806
rect 24332 5742 24334 5794
rect 24386 5742 24388 5794
rect 24332 5460 24388 5742
rect 24332 5404 25060 5460
rect 25004 5346 25060 5404
rect 25004 5294 25006 5346
rect 25058 5294 25060 5346
rect 25004 5282 25060 5294
rect 25340 5348 25396 5358
rect 25340 5346 25508 5348
rect 25340 5294 25342 5346
rect 25394 5294 25508 5346
rect 25340 5292 25508 5294
rect 25340 5282 25396 5292
rect 22988 5070 22990 5122
rect 23042 5070 23044 5122
rect 22540 5058 22596 5068
rect 22764 5058 22820 5068
rect 21420 4900 21476 4910
rect 21420 4806 21476 4844
rect 20748 4398 20750 4450
rect 20802 4398 20804 4450
rect 20748 4386 20804 4398
rect 19964 4340 20020 4350
rect 19628 4338 20020 4340
rect 19628 4286 19630 4338
rect 19682 4286 19966 4338
rect 20018 4286 20020 4338
rect 19628 4284 20020 4286
rect 19628 4274 19684 4284
rect 19964 4274 20020 4284
rect 22876 4228 22932 4238
rect 22988 4228 23044 5070
rect 22876 4226 23044 4228
rect 22876 4174 22878 4226
rect 22930 4174 23044 4226
rect 22876 4172 23044 4174
rect 23548 5236 23604 5246
rect 22876 4162 22932 4172
rect 18396 3602 18452 3612
rect 11900 3554 11956 3566
rect 11900 3502 11902 3554
rect 11954 3502 11956 3554
rect 11900 3444 11956 3502
rect 11900 3378 11956 3388
rect 12460 3444 12516 3454
rect 12460 3350 12516 3388
rect 23548 3444 23604 5180
rect 25340 5124 25396 5134
rect 25340 5030 25396 5068
rect 25340 4452 25396 4462
rect 25116 4450 25396 4452
rect 25116 4398 25342 4450
rect 25394 4398 25396 4450
rect 25116 4396 25396 4398
rect 24668 3556 24724 3566
rect 24668 3462 24724 3500
rect 23548 3378 23604 3388
rect 16156 3332 16212 3342
rect 16156 800 16212 3276
rect 16940 3332 16996 3342
rect 20860 3332 20916 3342
rect 16940 3238 16996 3276
rect 20636 3330 20916 3332
rect 20636 3278 20862 3330
rect 20914 3278 20916 3330
rect 20636 3276 20916 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20636 800 20692 3276
rect 20860 3266 20916 3276
rect 25116 800 25172 4396
rect 25340 4386 25396 4396
rect 25340 3668 25396 3678
rect 25452 3668 25508 5292
rect 25788 5124 25844 5134
rect 25788 5030 25844 5068
rect 26908 5124 26964 6636
rect 27020 6690 27076 6972
rect 27020 6638 27022 6690
rect 27074 6638 27076 6690
rect 27020 6626 27076 6638
rect 26908 5058 26964 5068
rect 27244 5908 27300 5918
rect 25340 3666 25508 3668
rect 25340 3614 25342 3666
rect 25394 3614 25508 3666
rect 25340 3612 25508 3614
rect 27244 3668 27300 5852
rect 27356 5906 27412 9548
rect 29036 9044 29092 15484
rect 29148 15314 29204 15326
rect 29148 15262 29150 15314
rect 29202 15262 29204 15314
rect 29148 15148 29204 15262
rect 29596 15316 29652 15326
rect 29596 15222 29652 15260
rect 29148 15092 29428 15148
rect 29372 14642 29428 15092
rect 29372 14590 29374 14642
rect 29426 14590 29428 14642
rect 29372 13300 29428 14590
rect 29484 14868 29540 14878
rect 29484 14308 29540 14812
rect 29484 13634 29540 14252
rect 29484 13582 29486 13634
rect 29538 13582 29540 13634
rect 29484 13570 29540 13582
rect 30156 14644 30212 14654
rect 29372 13234 29428 13244
rect 30156 13188 30212 14588
rect 30156 13122 30212 13132
rect 30268 12404 30324 17052
rect 30380 15202 30436 15214
rect 30380 15150 30382 15202
rect 30434 15150 30436 15202
rect 30380 14308 30436 15150
rect 30716 14308 30772 14318
rect 30380 14252 30716 14308
rect 30716 14242 30772 14252
rect 30268 12338 30324 12348
rect 30716 12962 30772 12974
rect 30716 12910 30718 12962
rect 30770 12910 30772 12962
rect 30716 12068 30772 12910
rect 30716 12002 30772 12012
rect 29484 11620 29540 11630
rect 29260 11396 29316 11406
rect 29260 11302 29316 11340
rect 29484 11396 29540 11564
rect 29484 11394 29764 11396
rect 29484 11342 29486 11394
rect 29538 11342 29764 11394
rect 29484 11340 29764 11342
rect 29484 11330 29540 11340
rect 29148 11282 29204 11294
rect 29148 11230 29150 11282
rect 29202 11230 29204 11282
rect 29148 9828 29204 11230
rect 29708 10498 29764 11340
rect 30380 10948 30436 10958
rect 30156 10836 30212 10846
rect 30380 10836 30436 10892
rect 29708 10446 29710 10498
rect 29762 10446 29764 10498
rect 29708 10434 29764 10446
rect 29932 10612 29988 10622
rect 29148 9714 29204 9772
rect 29484 10164 29540 10174
rect 29484 9940 29540 10108
rect 29932 9940 29988 10556
rect 30156 10610 30212 10780
rect 30156 10558 30158 10610
rect 30210 10558 30212 10610
rect 30156 10546 30212 10558
rect 30268 10834 30436 10836
rect 30268 10782 30382 10834
rect 30434 10782 30436 10834
rect 30268 10780 30436 10782
rect 30268 10164 30324 10780
rect 30380 10770 30436 10780
rect 30828 10836 30884 19852
rect 30940 19842 30996 19852
rect 31052 14868 31108 20524
rect 31276 18900 31332 25004
rect 31836 24948 31892 26852
rect 32172 26178 32228 26190
rect 32172 26126 32174 26178
rect 32226 26126 32228 26178
rect 32172 25732 32228 26126
rect 32172 25666 32228 25676
rect 31948 25620 32004 25630
rect 31948 25526 32004 25564
rect 31612 24892 31892 24948
rect 31612 23378 31668 24892
rect 32060 24836 32116 24846
rect 32060 24050 32116 24780
rect 32396 24836 32452 32732
rect 33292 32676 33348 34188
rect 33516 33908 33572 34300
rect 33628 34914 33684 34926
rect 33628 34862 33630 34914
rect 33682 34862 33684 34914
rect 33628 34354 33684 34862
rect 33964 34916 34020 35646
rect 34076 35364 34132 35758
rect 34300 35700 34356 35710
rect 34300 35698 34468 35700
rect 34300 35646 34302 35698
rect 34354 35646 34468 35698
rect 34300 35644 34468 35646
rect 34300 35634 34356 35644
rect 34412 35474 34468 35644
rect 34412 35422 34414 35474
rect 34466 35422 34468 35474
rect 34412 35410 34468 35422
rect 34636 35588 34692 35598
rect 34076 35298 34132 35308
rect 34636 35364 34692 35532
rect 34636 35298 34692 35308
rect 34748 35028 34804 42478
rect 34860 42978 34916 42990
rect 34860 42926 34862 42978
rect 34914 42926 34916 42978
rect 34860 42196 34916 42926
rect 34972 42644 35028 47012
rect 36988 46900 37044 47294
rect 37660 47346 37716 47358
rect 37660 47294 37662 47346
rect 37714 47294 37716 47346
rect 37324 47236 37380 47246
rect 37324 47142 37380 47180
rect 37100 46900 37156 46910
rect 36988 46898 37156 46900
rect 36988 46846 37102 46898
rect 37154 46846 37156 46898
rect 36988 46844 37156 46846
rect 37100 46834 37156 46844
rect 36428 46674 36484 46686
rect 36428 46622 36430 46674
rect 36482 46622 36484 46674
rect 36204 46564 36260 46574
rect 36428 46564 36484 46622
rect 36876 46676 36932 46686
rect 37436 46676 37492 46686
rect 36876 46582 36932 46620
rect 37324 46674 37492 46676
rect 37324 46622 37438 46674
rect 37490 46622 37492 46674
rect 37324 46620 37492 46622
rect 36204 46562 36484 46564
rect 36204 46510 36206 46562
rect 36258 46510 36484 46562
rect 36204 46508 36484 46510
rect 36988 46562 37044 46574
rect 36988 46510 36990 46562
rect 37042 46510 37044 46562
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35084 45778 35140 45790
rect 35084 45726 35086 45778
rect 35138 45726 35140 45778
rect 35084 45668 35140 45726
rect 35980 45780 36036 45790
rect 35084 45612 35364 45668
rect 35308 45108 35364 45612
rect 35308 45042 35364 45052
rect 35644 44994 35700 45006
rect 35644 44942 35646 44994
rect 35698 44942 35700 44994
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35532 44548 35588 44558
rect 35532 44454 35588 44492
rect 35084 44436 35140 44446
rect 35084 44342 35140 44380
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35084 42644 35140 42654
rect 34972 42588 35084 42644
rect 35084 42578 35140 42588
rect 34972 42196 35028 42206
rect 34860 42194 35028 42196
rect 34860 42142 34974 42194
rect 35026 42142 35028 42194
rect 34860 42140 35028 42142
rect 34972 42130 35028 42140
rect 35084 42084 35140 42094
rect 35084 41990 35140 42028
rect 34972 41748 35028 41758
rect 34972 41654 35028 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35644 40404 35700 44942
rect 35756 44212 35812 44222
rect 35756 44118 35812 44156
rect 35980 43428 36036 45724
rect 36092 45108 36148 45118
rect 36092 44322 36148 45052
rect 36092 44270 36094 44322
rect 36146 44270 36148 44322
rect 36092 43988 36148 44270
rect 36092 43922 36148 43932
rect 35980 43334 36036 43372
rect 36204 43204 36260 46508
rect 36428 46228 36484 46238
rect 36316 44322 36372 44334
rect 36316 44270 36318 44322
rect 36370 44270 36372 44322
rect 36316 43764 36372 44270
rect 36428 44098 36484 46172
rect 36988 45890 37044 46510
rect 36988 45838 36990 45890
rect 37042 45838 37044 45890
rect 36988 45826 37044 45838
rect 37212 45780 37268 45790
rect 37100 45778 37268 45780
rect 37100 45726 37214 45778
rect 37266 45726 37268 45778
rect 37100 45724 37268 45726
rect 37100 45108 37156 45724
rect 37212 45714 37268 45724
rect 37324 45780 37380 46620
rect 37436 46610 37492 46620
rect 37660 46228 37716 47294
rect 37772 47348 37828 47358
rect 37884 47348 37940 48860
rect 39004 48466 39060 49756
rect 39564 49746 39620 49756
rect 39788 49810 39844 49980
rect 41020 49970 41076 49982
rect 41132 49924 41188 49934
rect 41132 49830 41188 49868
rect 39788 49758 39790 49810
rect 39842 49758 39844 49810
rect 39788 48916 39844 49758
rect 40012 49810 40068 49822
rect 40012 49758 40014 49810
rect 40066 49758 40068 49810
rect 39900 49700 39956 49710
rect 39900 49606 39956 49644
rect 39788 48850 39844 48860
rect 39004 48414 39006 48466
rect 39058 48414 39060 48466
rect 39004 48402 39060 48414
rect 39228 48242 39284 48254
rect 39228 48190 39230 48242
rect 39282 48190 39284 48242
rect 39228 47684 39284 48190
rect 39228 47618 39284 47628
rect 39228 47458 39284 47470
rect 40012 47460 40068 49758
rect 39228 47406 39230 47458
rect 39282 47406 39284 47458
rect 38332 47348 38388 47358
rect 37772 47346 38500 47348
rect 37772 47294 37774 47346
rect 37826 47294 38334 47346
rect 38386 47294 38500 47346
rect 37772 47292 38500 47294
rect 37772 47282 37828 47292
rect 38332 47282 38388 47292
rect 38220 46564 38276 46574
rect 37548 46172 37660 46228
rect 37548 45890 37604 46172
rect 37660 46162 37716 46172
rect 38108 46562 38276 46564
rect 38108 46510 38222 46562
rect 38274 46510 38276 46562
rect 38108 46508 38276 46510
rect 37996 46004 38052 46014
rect 37548 45838 37550 45890
rect 37602 45838 37604 45890
rect 37548 45826 37604 45838
rect 37884 46002 38052 46004
rect 37884 45950 37998 46002
rect 38050 45950 38052 46002
rect 37884 45948 38052 45950
rect 37324 45714 37380 45724
rect 37884 45780 37940 45948
rect 37996 45938 38052 45948
rect 38108 45780 38164 46508
rect 38220 46498 38276 46508
rect 37884 45714 37940 45724
rect 37996 45724 38164 45780
rect 37436 45666 37492 45678
rect 37436 45614 37438 45666
rect 37490 45614 37492 45666
rect 37436 45556 37492 45614
rect 37996 45556 38052 45724
rect 37436 45500 38052 45556
rect 38332 45218 38388 45230
rect 38332 45166 38334 45218
rect 38386 45166 38388 45218
rect 37100 44436 37156 45052
rect 37212 45106 37268 45118
rect 37212 45054 37214 45106
rect 37266 45054 37268 45106
rect 37212 44996 37268 45054
rect 38220 45108 38276 45118
rect 38220 45014 38276 45052
rect 37212 44930 37268 44940
rect 37100 44370 37156 44380
rect 36428 44046 36430 44098
rect 36482 44046 36484 44098
rect 36428 44034 36484 44046
rect 37772 44212 37828 44222
rect 36316 43698 36372 43708
rect 37772 43538 37828 44156
rect 38220 44212 38276 44222
rect 38332 44212 38388 45166
rect 38444 44546 38500 47292
rect 39228 47236 39284 47406
rect 39452 47404 40068 47460
rect 39452 47346 39508 47404
rect 39452 47294 39454 47346
rect 39506 47294 39508 47346
rect 39452 47282 39508 47294
rect 38892 46340 38948 46350
rect 38892 45218 38948 46284
rect 38892 45166 38894 45218
rect 38946 45166 38948 45218
rect 38892 45154 38948 45166
rect 38444 44494 38446 44546
rect 38498 44494 38500 44546
rect 38444 44482 38500 44494
rect 38780 45108 38836 45118
rect 38780 44548 38836 45052
rect 38892 44548 38948 44558
rect 38780 44546 38948 44548
rect 38780 44494 38894 44546
rect 38946 44494 38948 44546
rect 38780 44492 38948 44494
rect 38892 44482 38948 44492
rect 38556 44324 38612 44334
rect 38556 44230 38612 44268
rect 39004 44324 39060 44334
rect 39004 44230 39060 44268
rect 38220 44210 38388 44212
rect 38220 44158 38222 44210
rect 38274 44158 38388 44210
rect 38220 44156 38388 44158
rect 37884 43876 37940 43886
rect 38220 43876 38276 44156
rect 37940 43820 38276 43876
rect 38780 43988 38836 43998
rect 37884 43650 37940 43820
rect 37884 43598 37886 43650
rect 37938 43598 37940 43650
rect 37884 43586 37940 43598
rect 37772 43486 37774 43538
rect 37826 43486 37828 43538
rect 37772 43474 37828 43486
rect 38780 43538 38836 43932
rect 39228 43762 39284 47180
rect 40012 47012 40068 47404
rect 40236 49810 40292 49822
rect 40236 49758 40238 49810
rect 40290 49758 40292 49810
rect 40236 47460 40292 49758
rect 40908 49700 40964 49710
rect 40908 49606 40964 49644
rect 40236 47394 40292 47404
rect 41132 48916 41188 48926
rect 40012 46946 40068 46956
rect 39900 46676 39956 46686
rect 39452 44994 39508 45006
rect 39452 44942 39454 44994
rect 39506 44942 39508 44994
rect 39452 44434 39508 44942
rect 39452 44382 39454 44434
rect 39506 44382 39508 44434
rect 39452 44324 39508 44382
rect 39508 44268 39620 44324
rect 39452 44258 39508 44268
rect 39228 43710 39230 43762
rect 39282 43710 39284 43762
rect 39228 43698 39284 43710
rect 39452 43764 39508 43774
rect 39452 43650 39508 43708
rect 39452 43598 39454 43650
rect 39506 43598 39508 43650
rect 39452 43586 39508 43598
rect 38780 43486 38782 43538
rect 38834 43486 38836 43538
rect 38780 43474 38836 43486
rect 36092 43148 36260 43204
rect 35868 42642 35924 42654
rect 35868 42590 35870 42642
rect 35922 42590 35924 42642
rect 35868 42532 35924 42590
rect 35980 42644 36036 42654
rect 35980 42550 36036 42588
rect 35868 42084 35924 42476
rect 36092 42308 36148 43148
rect 38556 42756 38612 42766
rect 38556 42662 38612 42700
rect 35868 42018 35924 42028
rect 35980 42252 36148 42308
rect 36204 42530 36260 42542
rect 36204 42478 36206 42530
rect 36258 42478 36260 42530
rect 35868 40404 35924 40414
rect 35532 40402 35924 40404
rect 35532 40350 35870 40402
rect 35922 40350 35924 40402
rect 35532 40348 35924 40350
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35420 38836 35476 38846
rect 35532 38836 35588 40348
rect 35868 40338 35924 40348
rect 35420 38834 35588 38836
rect 35420 38782 35422 38834
rect 35474 38782 35588 38834
rect 35420 38780 35588 38782
rect 35420 38770 35476 38780
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38164 35588 38780
rect 35980 38668 36036 42252
rect 36204 41188 36260 42478
rect 38220 42532 38276 42542
rect 38220 42438 38276 42476
rect 36204 41122 36260 41132
rect 36988 42308 37044 42318
rect 36652 40964 36708 40974
rect 36652 40514 36708 40908
rect 36652 40462 36654 40514
rect 36706 40462 36708 40514
rect 36652 40450 36708 40462
rect 36988 39844 37044 42252
rect 37100 41972 37156 41982
rect 37100 41186 37156 41916
rect 38108 41300 38164 41310
rect 37100 41134 37102 41186
rect 37154 41134 37156 41186
rect 37100 41076 37156 41134
rect 37212 41188 37268 41198
rect 37212 41094 37268 41132
rect 38108 41186 38164 41244
rect 38108 41134 38110 41186
rect 38162 41134 38164 41186
rect 38108 41122 38164 41134
rect 38556 41300 38612 41310
rect 37100 41010 37156 41020
rect 37548 41076 37604 41086
rect 37772 41076 37828 41086
rect 37548 41074 37828 41076
rect 37548 41022 37550 41074
rect 37602 41022 37774 41074
rect 37826 41022 37828 41074
rect 37548 41020 37828 41022
rect 37548 41010 37604 41020
rect 37772 41010 37828 41020
rect 37324 40964 37380 40974
rect 37324 40870 37380 40908
rect 37996 40962 38052 40974
rect 37996 40910 37998 40962
rect 38050 40910 38052 40962
rect 37996 40292 38052 40910
rect 38556 40740 38612 41244
rect 38556 40674 38612 40684
rect 39452 40962 39508 40974
rect 39452 40910 39454 40962
rect 39506 40910 39508 40962
rect 39452 40740 39508 40910
rect 39452 40674 39508 40684
rect 37996 40226 38052 40236
rect 38780 40292 38836 40302
rect 36988 39778 37044 39788
rect 38780 39172 38836 40236
rect 38780 39106 38836 39116
rect 39228 40290 39284 40302
rect 39228 40238 39230 40290
rect 39282 40238 39284 40290
rect 38108 38836 38164 38846
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35420 35700 35476 35710
rect 35532 35700 35588 38108
rect 35868 38612 36036 38668
rect 36092 38722 36148 38734
rect 36092 38670 36094 38722
rect 36146 38670 36148 38722
rect 36092 38668 36148 38670
rect 37212 38724 37268 38734
rect 36092 38612 36260 38668
rect 35420 35698 35532 35700
rect 35420 35646 35422 35698
rect 35474 35646 35532 35698
rect 35420 35644 35532 35646
rect 35588 35644 35700 35700
rect 35420 35634 35476 35644
rect 35532 35606 35588 35644
rect 34636 34972 34804 35028
rect 34860 35474 34916 35486
rect 35196 35476 35252 35486
rect 34860 35422 34862 35474
rect 34914 35422 34916 35474
rect 33964 34860 34132 34916
rect 33964 34692 34020 34702
rect 33628 34302 33630 34354
rect 33682 34302 33684 34354
rect 33628 34290 33684 34302
rect 33852 34690 34020 34692
rect 33852 34638 33966 34690
rect 34018 34638 34020 34690
rect 33852 34636 34020 34638
rect 33516 33842 33572 33852
rect 33852 33684 33908 34636
rect 33964 34626 34020 34636
rect 34076 34468 34132 34860
rect 34300 34804 34356 34814
rect 33964 34412 34132 34468
rect 34188 34690 34244 34702
rect 34188 34638 34190 34690
rect 34242 34638 34244 34690
rect 33964 34244 34020 34412
rect 34188 34356 34244 34638
rect 34188 34290 34244 34300
rect 34300 34354 34356 34748
rect 34524 34468 34580 34478
rect 34300 34302 34302 34354
rect 34354 34302 34356 34354
rect 34300 34290 34356 34302
rect 34412 34412 34524 34468
rect 33964 34150 34020 34188
rect 34076 34242 34132 34254
rect 34076 34190 34078 34242
rect 34130 34190 34132 34242
rect 34076 34132 34132 34190
rect 34412 34132 34468 34412
rect 34524 34402 34580 34412
rect 34076 34076 34468 34132
rect 34524 34132 34580 34142
rect 34524 34038 34580 34076
rect 34412 33908 34468 33918
rect 33852 33628 34132 33684
rect 33740 33572 33796 33582
rect 33516 33516 33740 33572
rect 33796 33516 33908 33572
rect 33516 32788 33572 33516
rect 33740 33506 33796 33516
rect 33852 33458 33908 33516
rect 33852 33406 33854 33458
rect 33906 33406 33908 33458
rect 33852 33394 33908 33406
rect 33964 33460 34020 33470
rect 33516 32694 33572 32732
rect 33404 32676 33460 32686
rect 33292 32674 33460 32676
rect 33292 32622 33406 32674
rect 33458 32622 33460 32674
rect 33292 32620 33460 32622
rect 33404 31666 33460 32620
rect 33740 32564 33796 32574
rect 33740 32562 33908 32564
rect 33740 32510 33742 32562
rect 33794 32510 33908 32562
rect 33740 32508 33908 32510
rect 33740 32498 33796 32508
rect 33852 31780 33908 32508
rect 33964 32562 34020 33404
rect 33964 32510 33966 32562
rect 34018 32510 34020 32562
rect 33964 32498 34020 32510
rect 33964 31780 34020 31790
rect 33852 31778 34020 31780
rect 33852 31726 33966 31778
rect 34018 31726 34020 31778
rect 33852 31724 34020 31726
rect 33964 31714 34020 31724
rect 33404 31614 33406 31666
rect 33458 31614 33460 31666
rect 33404 31602 33460 31614
rect 33068 31554 33124 31566
rect 33068 31502 33070 31554
rect 33122 31502 33124 31554
rect 33068 30884 33124 31502
rect 33628 31276 33908 31332
rect 33628 31106 33684 31276
rect 33628 31054 33630 31106
rect 33682 31054 33684 31106
rect 33628 31042 33684 31054
rect 33740 31106 33796 31118
rect 33740 31054 33742 31106
rect 33794 31054 33796 31106
rect 33068 30818 33124 30828
rect 32396 24770 32452 24780
rect 32508 29988 32564 29998
rect 32060 23998 32062 24050
rect 32114 23998 32116 24050
rect 32060 23986 32116 23998
rect 31612 23326 31614 23378
rect 31666 23326 31668 23378
rect 31612 23314 31668 23326
rect 31500 23156 31556 23166
rect 31388 23154 31556 23156
rect 31388 23102 31502 23154
rect 31554 23102 31556 23154
rect 31388 23100 31556 23102
rect 31388 19796 31444 23100
rect 31500 23090 31556 23100
rect 31500 22708 31556 22718
rect 31500 22484 31556 22652
rect 31500 22482 31892 22484
rect 31500 22430 31502 22482
rect 31554 22430 31892 22482
rect 31500 22428 31892 22430
rect 31500 22418 31556 22428
rect 31836 22370 31892 22428
rect 31836 22318 31838 22370
rect 31890 22318 31892 22370
rect 31836 22306 31892 22318
rect 32396 20916 32452 20926
rect 31836 20802 31892 20814
rect 31836 20750 31838 20802
rect 31890 20750 31892 20802
rect 31500 20580 31556 20590
rect 31500 20486 31556 20524
rect 31836 20356 31892 20750
rect 32060 20690 32116 20702
rect 32060 20638 32062 20690
rect 32114 20638 32116 20690
rect 32060 20580 32116 20638
rect 32060 20514 32116 20524
rect 31836 20300 32004 20356
rect 31836 20132 31892 20142
rect 31836 20038 31892 20076
rect 31948 20020 32004 20300
rect 32172 20020 32228 20030
rect 31948 19964 32172 20020
rect 32172 19926 32228 19964
rect 32396 20018 32452 20860
rect 32396 19966 32398 20018
rect 32450 19966 32452 20018
rect 32396 19954 32452 19966
rect 31388 19730 31444 19740
rect 32508 19460 32564 29932
rect 33740 29876 33796 31054
rect 33852 30996 33908 31276
rect 33964 31220 34020 31230
rect 34076 31220 34132 33628
rect 34412 33458 34468 33852
rect 34412 33406 34414 33458
rect 34466 33406 34468 33458
rect 34412 33394 34468 33406
rect 34636 32004 34692 34972
rect 34748 34804 34804 34814
rect 34860 34804 34916 35422
rect 35084 35420 35196 35476
rect 35084 35026 35140 35420
rect 35196 35410 35252 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34974 35086 35026
rect 35138 34974 35140 35026
rect 35084 34962 35140 34974
rect 34748 34802 34916 34804
rect 34748 34750 34750 34802
rect 34802 34750 34916 34802
rect 34748 34748 34916 34750
rect 35532 34804 35588 34814
rect 34748 34738 34804 34748
rect 35532 34710 35588 34748
rect 34972 34692 35028 34702
rect 34972 34690 35140 34692
rect 34972 34638 34974 34690
rect 35026 34638 35140 34690
rect 34972 34636 35140 34638
rect 34972 34626 35028 34636
rect 34860 34356 34916 34366
rect 34860 34242 34916 34300
rect 34860 34190 34862 34242
rect 34914 34190 34916 34242
rect 34636 31938 34692 31948
rect 34748 32450 34804 32462
rect 34748 32398 34750 32450
rect 34802 32398 34804 32450
rect 34636 31780 34692 31790
rect 34748 31780 34804 32398
rect 34636 31778 34804 31780
rect 34636 31726 34638 31778
rect 34690 31726 34804 31778
rect 34636 31724 34804 31726
rect 34636 31714 34692 31724
rect 34300 31556 34356 31566
rect 34524 31556 34580 31566
rect 34860 31556 34916 34190
rect 34300 31554 34468 31556
rect 34300 31502 34302 31554
rect 34354 31502 34468 31554
rect 34300 31500 34468 31502
rect 34300 31490 34356 31500
rect 33964 31218 34132 31220
rect 33964 31166 33966 31218
rect 34018 31166 34132 31218
rect 33964 31164 34132 31166
rect 34412 31220 34468 31500
rect 34524 31554 34916 31556
rect 34524 31502 34526 31554
rect 34578 31502 34916 31554
rect 34524 31500 34916 31502
rect 34972 34244 35028 34254
rect 34524 31490 34580 31500
rect 34524 31220 34580 31230
rect 34412 31218 34580 31220
rect 34412 31166 34526 31218
rect 34578 31166 34580 31218
rect 34412 31164 34580 31166
rect 33964 31154 34020 31164
rect 34524 31154 34580 31164
rect 34300 31108 34356 31118
rect 34972 31108 35028 34188
rect 34300 31014 34356 31052
rect 34636 31052 35028 31108
rect 34188 30996 34244 31006
rect 33852 30994 34244 30996
rect 33852 30942 34190 30994
rect 34242 30942 34244 30994
rect 33852 30940 34244 30942
rect 33740 29810 33796 29820
rect 34188 30212 34244 30940
rect 34076 29764 34132 29774
rect 33516 29540 33572 29550
rect 32732 28532 32788 28542
rect 32732 27412 32788 28476
rect 33516 28308 33572 29484
rect 33516 28242 33572 28252
rect 33628 28756 33684 28766
rect 32732 27186 32788 27356
rect 32732 27134 32734 27186
rect 32786 27134 32788 27186
rect 32732 27122 32788 27134
rect 33628 25284 33684 28700
rect 34076 28084 34132 29708
rect 34188 29650 34244 30156
rect 34636 29764 34692 31052
rect 34860 30882 34916 30894
rect 34860 30830 34862 30882
rect 34914 30830 34916 30882
rect 34860 29988 34916 30830
rect 35084 30436 35140 34636
rect 35196 34690 35252 34702
rect 35196 34638 35198 34690
rect 35250 34638 35252 34690
rect 35196 34356 35252 34638
rect 35196 34290 35252 34300
rect 35420 34468 35476 34478
rect 35420 34354 35476 34412
rect 35420 34302 35422 34354
rect 35474 34302 35476 34354
rect 35420 34290 35476 34302
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35644 33460 35700 35644
rect 35756 34690 35812 34702
rect 35756 34638 35758 34690
rect 35810 34638 35812 34690
rect 35756 34244 35812 34638
rect 35756 34178 35812 34188
rect 35868 34132 35924 38612
rect 35980 38500 36036 38510
rect 35980 38162 36036 38444
rect 35980 38110 35982 38162
rect 36034 38110 36036 38162
rect 35980 35140 36036 38110
rect 36092 35586 36148 35598
rect 36092 35534 36094 35586
rect 36146 35534 36148 35586
rect 36092 35476 36148 35534
rect 36092 35410 36148 35420
rect 35980 35074 36036 35084
rect 36092 35140 36148 35150
rect 36204 35140 36260 38612
rect 37100 38164 37156 38174
rect 37100 38070 37156 38108
rect 36092 35138 36260 35140
rect 36092 35086 36094 35138
rect 36146 35086 36260 35138
rect 36092 35084 36260 35086
rect 36092 35074 36148 35084
rect 35980 34690 36036 34702
rect 35980 34638 35982 34690
rect 36034 34638 36036 34690
rect 35980 34356 36036 34638
rect 37212 34468 37268 38668
rect 38108 37938 38164 38780
rect 38220 38724 38276 38762
rect 38892 38724 38948 38734
rect 39228 38724 39284 40238
rect 38220 38658 38276 38668
rect 38556 38722 39284 38724
rect 38556 38670 38894 38722
rect 38946 38670 39284 38722
rect 38556 38668 39284 38670
rect 39340 39172 39396 39182
rect 38556 38164 38612 38668
rect 38892 38658 38948 38668
rect 38556 38098 38612 38108
rect 39228 38162 39284 38174
rect 39228 38110 39230 38162
rect 39282 38110 39284 38162
rect 38108 37886 38110 37938
rect 38162 37886 38164 37938
rect 38108 37874 38164 37886
rect 37772 37826 37828 37838
rect 37772 37774 37774 37826
rect 37826 37774 37828 37826
rect 37436 37156 37492 37166
rect 37772 37156 37828 37774
rect 37212 34402 37268 34412
rect 37324 37154 37828 37156
rect 37324 37102 37438 37154
rect 37490 37102 37828 37154
rect 37324 37100 37828 37102
rect 35980 34290 36036 34300
rect 35644 33394 35700 33404
rect 35756 34020 35812 34030
rect 35868 34020 35924 34076
rect 35756 34018 35924 34020
rect 35756 33966 35758 34018
rect 35810 33966 35924 34018
rect 35756 33964 35924 33966
rect 35644 32340 35700 32350
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 31556 35588 31566
rect 35308 31108 35364 31118
rect 35308 31014 35364 31052
rect 35532 31108 35588 31500
rect 35532 31042 35588 31052
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30380 35252 30436
rect 34860 29922 34916 29932
rect 34188 29598 34190 29650
rect 34242 29598 34244 29650
rect 34188 29586 34244 29598
rect 34412 29708 34692 29764
rect 34300 29428 34356 29438
rect 34300 28754 34356 29372
rect 34300 28702 34302 28754
rect 34354 28702 34356 28754
rect 34300 28690 34356 28702
rect 34188 28084 34244 28094
rect 34076 28082 34244 28084
rect 34076 28030 34190 28082
rect 34242 28030 34244 28082
rect 34076 28028 34244 28030
rect 33628 25218 33684 25228
rect 33964 27860 34020 27870
rect 32620 24612 32676 24622
rect 32620 22482 32676 24556
rect 32620 22430 32622 22482
rect 32674 22430 32676 22482
rect 32620 22418 32676 22430
rect 32396 19404 32564 19460
rect 32732 21364 32788 21374
rect 31276 18834 31332 18844
rect 31836 18900 31892 18910
rect 31500 18676 31556 18686
rect 31388 18620 31500 18676
rect 31388 18562 31444 18620
rect 31500 18610 31556 18620
rect 31388 18510 31390 18562
rect 31442 18510 31444 18562
rect 31388 18498 31444 18510
rect 31724 18562 31780 18574
rect 31724 18510 31726 18562
rect 31778 18510 31780 18562
rect 31500 18452 31556 18462
rect 31500 18358 31556 18396
rect 31612 18340 31668 18350
rect 31612 18246 31668 18284
rect 31724 17892 31780 18510
rect 31836 18004 31892 18844
rect 32396 18674 32452 19404
rect 32732 19348 32788 21308
rect 33964 21028 34020 27804
rect 33964 20962 34020 20972
rect 32956 20916 33012 20926
rect 32956 20822 33012 20860
rect 33516 20802 33572 20814
rect 33516 20750 33518 20802
rect 33570 20750 33572 20802
rect 33516 20580 33572 20750
rect 33516 20514 33572 20524
rect 33180 20132 33236 20142
rect 33068 20020 33124 20030
rect 33068 19906 33124 19964
rect 33068 19854 33070 19906
rect 33122 19854 33124 19906
rect 33068 19842 33124 19854
rect 32732 19282 32788 19292
rect 32844 19684 32900 19694
rect 33180 19684 33236 20076
rect 32900 19628 33236 19684
rect 33404 19794 33460 19806
rect 33404 19742 33406 19794
rect 33458 19742 33460 19794
rect 32844 19346 32900 19628
rect 32844 19294 32846 19346
rect 32898 19294 32900 19346
rect 32844 19282 32900 19294
rect 32396 18622 32398 18674
rect 32450 18622 32452 18674
rect 31948 18564 32004 18574
rect 31948 18470 32004 18508
rect 32172 18452 32228 18462
rect 32172 18358 32228 18396
rect 31836 17938 31892 17948
rect 31724 17826 31780 17836
rect 32396 17668 32452 18622
rect 32508 19236 32564 19246
rect 32508 18564 32564 19180
rect 33404 19124 33460 19742
rect 33628 19236 33684 19246
rect 33628 19142 33684 19180
rect 33404 19058 33460 19068
rect 33740 19010 33796 19022
rect 33740 18958 33742 19010
rect 33794 18958 33796 19010
rect 33740 18900 33796 18958
rect 33740 18834 33796 18844
rect 33964 19010 34020 19022
rect 33964 18958 33966 19010
rect 34018 18958 34020 19010
rect 32508 18470 32564 18508
rect 33180 18450 33236 18462
rect 33180 18398 33182 18450
rect 33234 18398 33236 18450
rect 32620 17892 32676 17902
rect 32620 17798 32676 17836
rect 33180 17780 33236 18398
rect 33852 18340 33908 18350
rect 33180 17714 33236 17724
rect 33628 18338 33908 18340
rect 33628 18286 33854 18338
rect 33906 18286 33908 18338
rect 33628 18284 33908 18286
rect 33628 17778 33684 18284
rect 33852 18274 33908 18284
rect 33628 17726 33630 17778
rect 33682 17726 33684 17778
rect 33628 17714 33684 17726
rect 32396 17602 32452 17612
rect 33068 17668 33124 17678
rect 32732 17554 32788 17566
rect 32732 17502 32734 17554
rect 32786 17502 32788 17554
rect 32172 17442 32228 17454
rect 32172 17390 32174 17442
rect 32226 17390 32228 17442
rect 32172 17220 32228 17390
rect 32732 17220 32788 17502
rect 33068 17556 33124 17612
rect 33964 17666 34020 18958
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 33964 17602 34020 17614
rect 34076 18676 34132 28028
rect 34188 28018 34244 28028
rect 34412 27636 34468 29708
rect 35084 29652 35140 29662
rect 34524 29540 34580 29550
rect 34972 29540 35028 29550
rect 34524 29538 34916 29540
rect 34524 29486 34526 29538
rect 34578 29486 34916 29538
rect 34524 29484 34916 29486
rect 34524 29474 34580 29484
rect 34860 29426 34916 29484
rect 34972 29446 35028 29484
rect 34860 29374 34862 29426
rect 34914 29374 34916 29426
rect 34524 28196 34580 28206
rect 34524 28082 34580 28140
rect 34524 28030 34526 28082
rect 34578 28030 34580 28082
rect 34524 28018 34580 28030
rect 34860 27970 34916 29374
rect 34972 28756 35028 28766
rect 35084 28756 35140 29596
rect 35196 29650 35252 30380
rect 35644 29988 35700 32284
rect 35644 29922 35700 29932
rect 35196 29598 35198 29650
rect 35250 29598 35252 29650
rect 35196 29586 35252 29598
rect 35532 29540 35588 29550
rect 35532 29446 35588 29484
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35028 28700 35140 28756
rect 34972 28662 35028 28700
rect 35196 28196 35252 28206
rect 35084 28140 35196 28196
rect 34972 28084 35028 28094
rect 34972 27990 35028 28028
rect 34860 27918 34862 27970
rect 34914 27918 34916 27970
rect 34748 27860 34804 27870
rect 34860 27860 34916 27918
rect 34804 27804 34916 27860
rect 34748 27794 34804 27804
rect 34972 27636 35028 27646
rect 34412 27634 35028 27636
rect 34412 27582 34974 27634
rect 35026 27582 35028 27634
rect 34412 27580 35028 27582
rect 34972 27570 35028 27580
rect 34188 27412 34244 27422
rect 34188 25618 34244 27356
rect 34524 27076 34580 27086
rect 34524 26982 34580 27020
rect 35084 27074 35140 28140
rect 35196 28130 35252 28140
rect 35532 28196 35588 28206
rect 35756 28196 35812 33964
rect 37100 33236 37156 33246
rect 36988 32788 37044 32798
rect 36988 32694 37044 32732
rect 37100 31780 37156 33180
rect 37212 33124 37268 33134
rect 37212 33030 37268 33068
rect 36988 31724 37156 31780
rect 37212 32002 37268 32014
rect 37212 31950 37214 32002
rect 37266 31950 37268 32002
rect 36876 29988 36932 29998
rect 35868 29876 35924 29886
rect 35868 28756 35924 29820
rect 35980 29652 36036 29662
rect 35980 29426 36036 29596
rect 35980 29374 35982 29426
rect 36034 29374 36036 29426
rect 35980 29362 36036 29374
rect 36652 29314 36708 29326
rect 36652 29262 36654 29314
rect 36706 29262 36708 29314
rect 36652 28756 36708 29262
rect 35868 28754 36372 28756
rect 35868 28702 35870 28754
rect 35922 28702 36372 28754
rect 35868 28700 36372 28702
rect 35868 28690 35924 28700
rect 36204 28530 36260 28542
rect 36204 28478 36206 28530
rect 36258 28478 36260 28530
rect 35588 28140 35924 28196
rect 35532 28082 35588 28140
rect 35532 28030 35534 28082
rect 35586 28030 35588 28082
rect 35532 28018 35588 28030
rect 35644 27860 35700 27870
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35084 27022 35086 27074
rect 35138 27022 35140 27074
rect 35084 27010 35140 27022
rect 35644 27076 35700 27804
rect 34188 25566 34190 25618
rect 34242 25566 34244 25618
rect 34188 25554 34244 25566
rect 34412 26964 34468 26974
rect 34412 24834 34468 26908
rect 34860 26964 34916 27002
rect 35644 26982 35700 27020
rect 35868 27076 35924 28140
rect 35980 28084 36036 28094
rect 35980 27524 36036 28028
rect 36204 27748 36260 28478
rect 36316 28532 36372 28700
rect 36652 28690 36708 28700
rect 36540 28644 36596 28654
rect 36876 28644 36932 29932
rect 36988 28756 37044 31724
rect 37100 31556 37156 31566
rect 37212 31556 37268 31950
rect 37324 31668 37380 37100
rect 37436 37090 37492 37100
rect 39228 36932 39284 38110
rect 39228 36866 39284 36876
rect 39116 36484 39172 36494
rect 39116 36390 39172 36428
rect 39340 36482 39396 39116
rect 39564 38668 39620 44268
rect 39788 44210 39844 44222
rect 39788 44158 39790 44210
rect 39842 44158 39844 44210
rect 39788 44100 39844 44158
rect 39900 44210 39956 46620
rect 40348 46676 40404 46686
rect 40348 46562 40404 46620
rect 40348 46510 40350 46562
rect 40402 46510 40404 46562
rect 40348 46498 40404 46510
rect 39900 44158 39902 44210
rect 39954 44158 39956 44210
rect 39900 44146 39956 44158
rect 40012 45332 40068 45342
rect 41132 45332 41188 48860
rect 41580 46788 41636 46798
rect 41580 46694 41636 46732
rect 41244 46676 41300 46686
rect 41244 46582 41300 46620
rect 41244 45332 41300 45342
rect 41132 45330 41300 45332
rect 41132 45278 41246 45330
rect 41298 45278 41300 45330
rect 41132 45276 41300 45278
rect 39788 44034 39844 44044
rect 40012 43764 40068 45276
rect 41244 45266 41300 45276
rect 41132 45106 41188 45118
rect 41132 45054 41134 45106
rect 41186 45054 41188 45106
rect 40684 44324 40740 44334
rect 40684 44210 40740 44268
rect 41132 44324 41188 45054
rect 41132 44258 41188 44268
rect 41244 44882 41300 44894
rect 41244 44830 41246 44882
rect 41298 44830 41300 44882
rect 40684 44158 40686 44210
rect 40738 44158 40740 44210
rect 40684 44146 40740 44158
rect 40012 43538 40068 43708
rect 40124 44098 40180 44110
rect 40124 44046 40126 44098
rect 40178 44046 40180 44098
rect 40124 43708 40180 44046
rect 40348 44100 40404 44110
rect 40124 43652 40292 43708
rect 40012 43486 40014 43538
rect 40066 43486 40068 43538
rect 39788 43428 39844 43438
rect 39844 43372 39956 43428
rect 39788 43334 39844 43372
rect 39900 42642 39956 43372
rect 40012 42754 40068 43486
rect 40012 42702 40014 42754
rect 40066 42702 40068 42754
rect 40012 42690 40068 42702
rect 39900 42590 39902 42642
rect 39954 42590 39956 42642
rect 39900 42578 39956 42590
rect 39676 42530 39732 42542
rect 39676 42478 39678 42530
rect 39730 42478 39732 42530
rect 39676 41186 39732 42478
rect 40236 42084 40292 43652
rect 40348 43314 40404 44044
rect 40348 43262 40350 43314
rect 40402 43262 40404 43314
rect 40348 42756 40404 43262
rect 41132 43426 41188 43438
rect 41132 43374 41134 43426
rect 41186 43374 41188 43426
rect 41132 42980 41188 43374
rect 41132 42914 41188 42924
rect 40348 42690 40404 42700
rect 40236 42028 40852 42084
rect 39676 41134 39678 41186
rect 39730 41134 39732 41186
rect 39676 40628 39732 41134
rect 40124 41300 40180 41310
rect 40124 41186 40180 41244
rect 40124 41134 40126 41186
rect 40178 41134 40180 41186
rect 40124 41122 40180 41134
rect 39676 40562 39732 40572
rect 40124 40628 40180 40638
rect 40124 38946 40180 40572
rect 40796 39284 40852 42028
rect 41244 42082 41300 44830
rect 41356 44322 41412 44334
rect 41356 44270 41358 44322
rect 41410 44270 41412 44322
rect 41356 43652 41412 44270
rect 41692 43708 41748 51212
rect 41916 51202 41972 51212
rect 48636 50706 48692 50718
rect 48636 50654 48638 50706
rect 48690 50654 48692 50706
rect 42700 50596 42756 50606
rect 42364 50484 42420 50494
rect 42364 50390 42420 50428
rect 42028 49924 42084 49934
rect 42364 49924 42420 49934
rect 42028 49810 42084 49868
rect 42028 49758 42030 49810
rect 42082 49758 42084 49810
rect 42028 48804 42084 49758
rect 42252 49868 42364 49924
rect 42252 49810 42308 49868
rect 42364 49858 42420 49868
rect 42252 49758 42254 49810
rect 42306 49758 42308 49810
rect 42252 49746 42308 49758
rect 42700 49810 42756 50540
rect 43036 50596 43092 50606
rect 43036 50502 43092 50540
rect 43372 50596 43428 50606
rect 42700 49758 42702 49810
rect 42754 49758 42756 49810
rect 42700 49746 42756 49758
rect 42364 49588 42420 49598
rect 42364 49586 42644 49588
rect 42364 49534 42366 49586
rect 42418 49534 42644 49586
rect 42364 49532 42644 49534
rect 42364 49522 42420 49532
rect 42252 48916 42308 48926
rect 42252 48822 42308 48860
rect 42028 48738 42084 48748
rect 42476 48804 42532 48814
rect 42476 48710 42532 48748
rect 42588 48356 42644 49532
rect 42476 48300 42644 48356
rect 42700 49026 42756 49038
rect 42700 48974 42702 49026
rect 42754 48974 42756 49026
rect 42700 48916 42756 48974
rect 42364 47684 42420 47694
rect 42364 47460 42420 47628
rect 42476 47570 42532 48300
rect 42476 47518 42478 47570
rect 42530 47518 42532 47570
rect 42476 47506 42532 47518
rect 42140 47458 42420 47460
rect 42140 47406 42366 47458
rect 42418 47406 42420 47458
rect 42140 47404 42420 47406
rect 41804 47012 41860 47022
rect 41804 46898 41860 46956
rect 41804 46846 41806 46898
rect 41858 46846 41860 46898
rect 41804 46788 41860 46846
rect 42140 46898 42196 47404
rect 42364 47394 42420 47404
rect 42588 47460 42644 47470
rect 42588 47366 42644 47404
rect 42700 47124 42756 48860
rect 43148 47684 43204 47694
rect 42924 47458 42980 47470
rect 42924 47406 42926 47458
rect 42978 47406 42980 47458
rect 42812 47236 42868 47246
rect 42812 47142 42868 47180
rect 42140 46846 42142 46898
rect 42194 46846 42196 46898
rect 42140 46834 42196 46846
rect 42476 47068 42756 47124
rect 41804 46722 41860 46732
rect 42028 46674 42084 46686
rect 42028 46622 42030 46674
rect 42082 46622 42084 46674
rect 41916 46562 41972 46574
rect 41916 46510 41918 46562
rect 41970 46510 41972 46562
rect 41804 46452 41860 46462
rect 41916 46452 41972 46510
rect 42028 46564 42084 46622
rect 42028 46508 42420 46564
rect 41916 46396 42308 46452
rect 41804 45332 41860 46396
rect 41916 45332 41972 45342
rect 41804 45330 41972 45332
rect 41804 45278 41918 45330
rect 41970 45278 41972 45330
rect 41804 45276 41972 45278
rect 41916 45108 41972 45276
rect 42252 45218 42308 46396
rect 42252 45166 42254 45218
rect 42306 45166 42308 45218
rect 42252 45154 42308 45166
rect 42364 45778 42420 46508
rect 42364 45726 42366 45778
rect 42418 45726 42420 45778
rect 42364 45220 42420 45726
rect 42476 45668 42532 47068
rect 42924 47012 42980 47406
rect 42812 46956 42980 47012
rect 42588 46788 42644 46798
rect 42588 45890 42644 46732
rect 42700 46450 42756 46462
rect 42700 46398 42702 46450
rect 42754 46398 42756 46450
rect 42700 46002 42756 46398
rect 42700 45950 42702 46002
rect 42754 45950 42756 46002
rect 42700 45938 42756 45950
rect 42588 45838 42590 45890
rect 42642 45838 42644 45890
rect 42588 45826 42644 45838
rect 42812 45892 42868 46956
rect 42924 46786 42980 46798
rect 42924 46734 42926 46786
rect 42978 46734 42980 46786
rect 42924 46676 42980 46734
rect 42924 46610 42980 46620
rect 43036 46564 43092 46574
rect 43036 46470 43092 46508
rect 42812 45798 42868 45836
rect 43036 45892 43092 45902
rect 43148 45892 43204 47628
rect 43372 46676 43428 50540
rect 45724 50596 45780 50606
rect 45724 50502 45780 50540
rect 46508 50482 46564 50494
rect 46508 50430 46510 50482
rect 46562 50430 46564 50482
rect 43484 49924 43540 49934
rect 43484 49830 43540 49868
rect 46060 49812 46116 49822
rect 45612 49700 45668 49710
rect 45500 49698 45668 49700
rect 45500 49646 45614 49698
rect 45666 49646 45668 49698
rect 45500 49644 45668 49646
rect 45500 47460 45556 49644
rect 45612 49634 45668 49644
rect 46060 49028 46116 49756
rect 43372 46582 43428 46620
rect 45276 46676 45332 46686
rect 44156 46564 44212 46574
rect 44156 46470 44212 46508
rect 43036 45890 43204 45892
rect 43036 45838 43038 45890
rect 43090 45838 43204 45890
rect 43036 45836 43204 45838
rect 43036 45826 43092 45836
rect 42476 45612 42644 45668
rect 42364 45154 42420 45164
rect 42476 45218 42532 45230
rect 42476 45166 42478 45218
rect 42530 45166 42532 45218
rect 41692 43652 41860 43708
rect 41356 43586 41412 43596
rect 41468 43540 41524 43550
rect 41468 42980 41524 43484
rect 41468 42914 41524 42924
rect 41244 42030 41246 42082
rect 41298 42030 41300 42082
rect 41244 42018 41300 42030
rect 41020 41972 41076 41982
rect 41020 41878 41076 41916
rect 41692 41970 41748 41982
rect 41692 41918 41694 41970
rect 41746 41918 41748 41970
rect 41468 41860 41524 41870
rect 41132 41858 41524 41860
rect 41132 41806 41470 41858
rect 41522 41806 41524 41858
rect 41132 41804 41524 41806
rect 41132 41412 41188 41804
rect 41468 41794 41524 41804
rect 40908 41356 41188 41412
rect 40908 41298 40964 41356
rect 40908 41246 40910 41298
rect 40962 41246 40964 41298
rect 40908 41234 40964 41246
rect 40908 40628 40964 40638
rect 40908 40534 40964 40572
rect 41692 40626 41748 41918
rect 41692 40574 41694 40626
rect 41746 40574 41748 40626
rect 41692 40562 41748 40574
rect 41244 40514 41300 40526
rect 41244 40462 41246 40514
rect 41298 40462 41300 40514
rect 41244 40292 41300 40462
rect 41244 40226 41300 40236
rect 40796 39228 41300 39284
rect 41132 39058 41188 39070
rect 41132 39006 41134 39058
rect 41186 39006 41188 39058
rect 40124 38894 40126 38946
rect 40178 38894 40180 38946
rect 40124 38882 40180 38894
rect 40236 38946 40292 38958
rect 40236 38894 40238 38946
rect 40290 38894 40292 38946
rect 39564 38612 40068 38668
rect 39340 36430 39342 36482
rect 39394 36430 39396 36482
rect 39340 36418 39396 36430
rect 38332 36260 38388 36270
rect 38332 36166 38388 36204
rect 38780 36258 38836 36270
rect 38780 36206 38782 36258
rect 38834 36206 38836 36258
rect 38220 35588 38276 35598
rect 38276 35532 38500 35588
rect 38220 35494 38276 35532
rect 37884 35140 37940 35150
rect 37436 35028 37492 35038
rect 37492 34972 37604 35028
rect 37436 34962 37492 34972
rect 37548 33684 37604 34972
rect 37884 34356 37940 35084
rect 38444 35026 38500 35532
rect 38780 35252 38836 36206
rect 38892 36260 38948 36270
rect 38892 36166 38948 36204
rect 39004 36258 39060 36270
rect 39004 36206 39006 36258
rect 39058 36206 39060 36258
rect 38892 35700 38948 35710
rect 38892 35606 38948 35644
rect 38780 35186 38836 35196
rect 39004 35140 39060 36206
rect 39452 35700 39508 35710
rect 39004 35074 39060 35084
rect 39340 35644 39452 35700
rect 38444 34974 38446 35026
rect 38498 34974 38500 35026
rect 38444 34580 38500 34974
rect 38780 35028 38836 35038
rect 38444 34514 38500 34524
rect 38556 34692 38612 34702
rect 37884 34262 37940 34300
rect 38444 34356 38500 34366
rect 38556 34356 38612 34636
rect 38444 34354 38612 34356
rect 38444 34302 38446 34354
rect 38498 34302 38612 34354
rect 38444 34300 38612 34302
rect 38780 34692 38836 34972
rect 39228 35028 39284 35038
rect 38780 34356 38836 34636
rect 38444 34290 38500 34300
rect 38668 34244 38724 34254
rect 38668 34150 38724 34188
rect 38220 34132 38276 34142
rect 37436 33460 37492 33470
rect 37436 31780 37492 33404
rect 37548 32786 37604 33628
rect 37548 32734 37550 32786
rect 37602 32734 37604 32786
rect 37548 32722 37604 32734
rect 37996 34130 38276 34132
rect 37996 34078 38222 34130
rect 38274 34078 38276 34130
rect 37996 34076 38276 34078
rect 37772 32676 37828 32686
rect 37660 32564 37716 32574
rect 37548 32562 37716 32564
rect 37548 32510 37662 32562
rect 37714 32510 37716 32562
rect 37548 32508 37716 32510
rect 37548 32002 37604 32508
rect 37660 32498 37716 32508
rect 37772 32562 37828 32620
rect 37772 32510 37774 32562
rect 37826 32510 37828 32562
rect 37772 32498 37828 32510
rect 37884 32562 37940 32574
rect 37884 32510 37886 32562
rect 37938 32510 37940 32562
rect 37884 32452 37940 32510
rect 37884 32386 37940 32396
rect 37548 31950 37550 32002
rect 37602 31950 37604 32002
rect 37548 31938 37604 31950
rect 37660 31890 37716 31902
rect 37660 31838 37662 31890
rect 37714 31838 37716 31890
rect 37660 31780 37716 31838
rect 37436 31724 37716 31780
rect 37324 31612 37940 31668
rect 37100 31554 37268 31556
rect 37100 31502 37102 31554
rect 37154 31502 37268 31554
rect 37100 31500 37268 31502
rect 37100 29428 37156 31500
rect 37100 29362 37156 29372
rect 37324 28756 37380 28766
rect 36988 28700 37156 28756
rect 36540 28550 36596 28588
rect 36764 28588 37044 28644
rect 36316 28530 36484 28532
rect 36316 28478 36318 28530
rect 36370 28478 36484 28530
rect 36316 28476 36484 28478
rect 36316 28466 36372 28476
rect 36428 27860 36484 28476
rect 36764 28082 36820 28588
rect 36988 28530 37044 28588
rect 36988 28478 36990 28530
rect 37042 28478 37044 28530
rect 36988 28466 37044 28478
rect 37100 28308 37156 28700
rect 37212 28644 37268 28654
rect 37324 28644 37380 28700
rect 37436 28644 37492 28654
rect 37324 28642 37492 28644
rect 37324 28590 37438 28642
rect 37490 28590 37492 28642
rect 37324 28588 37492 28590
rect 37212 28550 37268 28588
rect 37436 28578 37492 28588
rect 37548 28644 37604 28654
rect 37772 28644 37828 28654
rect 37548 28642 37828 28644
rect 37548 28590 37550 28642
rect 37602 28590 37774 28642
rect 37826 28590 37828 28642
rect 37548 28588 37828 28590
rect 37548 28578 37604 28588
rect 37772 28578 37828 28588
rect 37884 28420 37940 31612
rect 36764 28030 36766 28082
rect 36818 28030 36820 28082
rect 36764 28018 36820 28030
rect 36988 28252 37156 28308
rect 37772 28364 37940 28420
rect 37996 28644 38052 34076
rect 38220 34066 38276 34076
rect 38556 34132 38612 34142
rect 38556 34038 38612 34076
rect 38444 33684 38500 33694
rect 38108 33124 38164 33134
rect 38108 32564 38164 33068
rect 38108 32562 38388 32564
rect 38108 32510 38110 32562
rect 38162 32510 38388 32562
rect 38108 32508 38388 32510
rect 38108 32498 38164 32508
rect 37996 28530 38052 28588
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 36428 27804 36708 27860
rect 36204 27692 36484 27748
rect 35980 27458 36036 27468
rect 34860 26898 34916 26908
rect 35868 26962 35924 27020
rect 35868 26910 35870 26962
rect 35922 26910 35924 26962
rect 35868 26898 35924 26910
rect 36092 27188 36148 27198
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34860 25732 34916 25742
rect 34748 25284 34804 25294
rect 34748 25190 34804 25228
rect 34412 24782 34414 24834
rect 34466 24782 34468 24834
rect 34412 23940 34468 24782
rect 34748 24836 34804 24846
rect 34860 24836 34916 25676
rect 35196 25730 35252 25742
rect 35196 25678 35198 25730
rect 35250 25678 35252 25730
rect 35084 25620 35140 25630
rect 34972 25172 35028 25182
rect 34972 24946 35028 25116
rect 34972 24894 34974 24946
rect 35026 24894 35028 24946
rect 34972 24882 35028 24894
rect 34748 24834 34916 24836
rect 34748 24782 34750 24834
rect 34802 24782 34916 24834
rect 34748 24780 34916 24782
rect 34524 24722 34580 24734
rect 34524 24670 34526 24722
rect 34578 24670 34580 24722
rect 34524 23940 34580 24670
rect 34636 24612 34692 24622
rect 34636 24518 34692 24556
rect 34636 23940 34692 23950
rect 34524 23938 34692 23940
rect 34524 23886 34638 23938
rect 34690 23886 34692 23938
rect 34524 23884 34692 23886
rect 34412 23874 34468 23884
rect 34636 23874 34692 23884
rect 34748 23716 34804 24780
rect 34972 24052 35028 24062
rect 34972 23938 35028 23996
rect 34972 23886 34974 23938
rect 35026 23886 35028 23938
rect 34972 23874 35028 23886
rect 34636 23660 34804 23716
rect 34860 23714 34916 23726
rect 34860 23662 34862 23714
rect 34914 23662 34916 23714
rect 34300 21474 34356 21486
rect 34300 21422 34302 21474
rect 34354 21422 34356 21474
rect 34300 21364 34356 21422
rect 34300 20132 34356 21308
rect 34300 20066 34356 20076
rect 34524 20578 34580 20590
rect 34524 20526 34526 20578
rect 34578 20526 34580 20578
rect 34524 19236 34580 20526
rect 34636 20020 34692 23660
rect 34748 22484 34804 22494
rect 34860 22484 34916 23662
rect 34748 22482 34916 22484
rect 34748 22430 34750 22482
rect 34802 22430 34916 22482
rect 34748 22428 34916 22430
rect 34748 21812 34804 22428
rect 34748 20580 34804 21756
rect 34860 21588 34916 21598
rect 34860 21494 34916 21532
rect 34860 20804 34916 20814
rect 35084 20804 35140 25564
rect 35196 25618 35252 25678
rect 35196 25566 35198 25618
rect 35250 25566 35252 25618
rect 35196 25554 35252 25566
rect 35532 25284 35588 25294
rect 35532 24724 35588 25228
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35308 21700 35364 21710
rect 35308 21606 35364 21644
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34860 20802 35140 20804
rect 34860 20750 34862 20802
rect 34914 20750 35140 20802
rect 34860 20748 35140 20750
rect 34860 20738 34916 20748
rect 34748 20524 35028 20580
rect 34748 20020 34804 20030
rect 34636 19964 34748 20020
rect 34748 19954 34804 19964
rect 34412 19180 34524 19236
rect 34300 19010 34356 19022
rect 34300 18958 34302 19010
rect 34354 18958 34356 19010
rect 34300 18900 34356 18958
rect 34300 18834 34356 18844
rect 33180 17556 33236 17566
rect 33068 17554 33236 17556
rect 33068 17502 33182 17554
rect 33234 17502 33236 17554
rect 33068 17500 33236 17502
rect 32172 17164 32732 17220
rect 32284 17106 32340 17164
rect 32732 17154 32788 17164
rect 33180 17332 33236 17500
rect 33852 17554 33908 17566
rect 33852 17502 33854 17554
rect 33906 17502 33908 17554
rect 33852 17444 33908 17502
rect 34076 17444 34132 18620
rect 34412 17666 34468 19180
rect 34524 19170 34580 19180
rect 34412 17614 34414 17666
rect 34466 17614 34468 17666
rect 34412 17602 34468 17614
rect 33852 17388 34132 17444
rect 34188 17444 34244 17454
rect 34188 17350 34244 17388
rect 32284 17054 32286 17106
rect 32338 17054 32340 17106
rect 32284 17042 32340 17054
rect 32060 15316 32116 15326
rect 31052 14802 31108 14812
rect 31164 14980 31220 14990
rect 31164 14644 31220 14924
rect 31164 14642 31556 14644
rect 31164 14590 31166 14642
rect 31218 14590 31556 14642
rect 31164 14588 31556 14590
rect 31164 14578 31220 14588
rect 31500 14530 31556 14588
rect 31500 14478 31502 14530
rect 31554 14478 31556 14530
rect 31500 14466 31556 14478
rect 31836 14530 31892 14542
rect 31836 14478 31838 14530
rect 31890 14478 31892 14530
rect 31500 14308 31556 14318
rect 31500 14214 31556 14252
rect 31836 13076 31892 14478
rect 32060 14530 32116 15260
rect 32508 15204 32564 15242
rect 32508 15138 32564 15148
rect 32060 14478 32062 14530
rect 32114 14478 32116 14530
rect 32060 14466 32116 14478
rect 32284 14420 32340 14430
rect 31836 13010 31892 13020
rect 32172 14418 32340 14420
rect 32172 14366 32286 14418
rect 32338 14366 32340 14418
rect 32172 14364 32340 14366
rect 31500 12852 31556 12862
rect 31500 12850 31892 12852
rect 31500 12798 31502 12850
rect 31554 12798 31892 12850
rect 31500 12796 31892 12798
rect 31500 12786 31556 12796
rect 31836 12402 31892 12796
rect 32172 12404 32228 14364
rect 32284 14354 32340 14364
rect 33180 13188 33236 17276
rect 34188 16884 34244 16894
rect 33404 15428 33460 15438
rect 33964 15428 34020 15438
rect 33404 15426 34020 15428
rect 33404 15374 33406 15426
rect 33458 15374 33966 15426
rect 34018 15374 34020 15426
rect 33404 15372 34020 15374
rect 33404 15204 33460 15372
rect 33964 15362 34020 15372
rect 33404 15138 33460 15148
rect 33516 15204 33572 15214
rect 33740 15204 33796 15214
rect 33516 15202 33740 15204
rect 33516 15150 33518 15202
rect 33570 15150 33740 15202
rect 33516 15148 33740 15150
rect 33516 15138 33572 15148
rect 33740 15138 33796 15148
rect 33180 13122 33236 13132
rect 33628 13074 33684 13086
rect 33628 13022 33630 13074
rect 33682 13022 33684 13074
rect 33628 12964 33684 13022
rect 33628 12898 33684 12908
rect 31836 12350 31838 12402
rect 31890 12350 31892 12402
rect 31836 12338 31892 12350
rect 31948 12348 32228 12404
rect 31724 11954 31780 11966
rect 31724 11902 31726 11954
rect 31778 11902 31780 11954
rect 31724 11506 31780 11902
rect 31948 11956 32004 12348
rect 32060 12178 32116 12190
rect 32060 12126 32062 12178
rect 32114 12126 32116 12178
rect 32060 12068 32116 12126
rect 33852 12180 33908 12190
rect 32060 12012 32564 12068
rect 31948 11900 32228 11956
rect 31724 11454 31726 11506
rect 31778 11454 31780 11506
rect 31724 11442 31780 11454
rect 30940 11396 30996 11406
rect 31164 11396 31220 11406
rect 30940 11394 31220 11396
rect 30940 11342 30942 11394
rect 30994 11342 31166 11394
rect 31218 11342 31220 11394
rect 30940 11340 31220 11342
rect 30940 11330 30996 11340
rect 30940 10836 30996 10846
rect 30884 10834 30996 10836
rect 30884 10782 30942 10834
rect 30994 10782 30996 10834
rect 30884 10780 30996 10782
rect 30828 10742 30884 10780
rect 30940 10770 30996 10780
rect 31164 10724 31220 11340
rect 31612 11396 31668 11406
rect 31612 11302 31668 11340
rect 31948 11396 32004 11406
rect 31164 10658 31220 10668
rect 31836 11170 31892 11182
rect 31836 11118 31838 11170
rect 31890 11118 31892 11170
rect 31836 10722 31892 11118
rect 31948 10834 32004 11340
rect 31948 10782 31950 10834
rect 32002 10782 32004 10834
rect 31948 10770 32004 10782
rect 32172 11394 32228 11900
rect 32508 11506 32564 12012
rect 32508 11454 32510 11506
rect 32562 11454 32564 11506
rect 32508 11442 32564 11454
rect 32172 11342 32174 11394
rect 32226 11342 32228 11394
rect 32172 10834 32228 11342
rect 32620 11396 32676 11406
rect 32620 11302 32676 11340
rect 32844 11394 32900 11406
rect 32844 11342 32846 11394
rect 32898 11342 32900 11394
rect 32844 11284 32900 11342
rect 32844 11218 32900 11228
rect 32396 11172 32452 11182
rect 32396 11078 32452 11116
rect 33404 11172 33460 11182
rect 32172 10782 32174 10834
rect 32226 10782 32228 10834
rect 32172 10770 32228 10782
rect 31836 10670 31838 10722
rect 31890 10670 31892 10722
rect 29484 9938 29988 9940
rect 29484 9886 29934 9938
rect 29986 9886 29988 9938
rect 29484 9884 29988 9886
rect 29484 9826 29540 9884
rect 29932 9874 29988 9884
rect 30044 10108 30324 10164
rect 29484 9774 29486 9826
rect 29538 9774 29540 9826
rect 29484 9762 29540 9774
rect 29148 9662 29150 9714
rect 29202 9662 29204 9714
rect 29148 9650 29204 9662
rect 29820 9268 29876 9278
rect 30044 9268 30100 10108
rect 31724 9268 31780 9278
rect 29820 9266 30100 9268
rect 29820 9214 29822 9266
rect 29874 9214 30100 9266
rect 29820 9212 30100 9214
rect 31612 9266 31780 9268
rect 31612 9214 31726 9266
rect 31778 9214 31780 9266
rect 31612 9212 31780 9214
rect 29820 9202 29876 9212
rect 29260 9044 29316 9054
rect 29036 9042 29316 9044
rect 29036 8990 29262 9042
rect 29314 8990 29316 9042
rect 29036 8988 29316 8990
rect 29036 8372 29092 8988
rect 29260 8978 29316 8988
rect 31052 9044 31108 9054
rect 31388 9044 31444 9054
rect 31052 9042 31444 9044
rect 31052 8990 31054 9042
rect 31106 8990 31390 9042
rect 31442 8990 31444 9042
rect 31052 8988 31444 8990
rect 31052 8978 31108 8988
rect 29036 8306 29092 8316
rect 30828 8258 30884 8270
rect 30828 8206 30830 8258
rect 30882 8206 30884 8258
rect 28700 8036 28756 8046
rect 28700 7586 28756 7980
rect 28700 7534 28702 7586
rect 28754 7534 28756 7586
rect 28700 7522 28756 7534
rect 29484 7474 29540 7486
rect 29484 7422 29486 7474
rect 29538 7422 29540 7474
rect 29484 7364 29540 7422
rect 29484 7298 29540 7308
rect 30828 7364 30884 8206
rect 31164 7700 31220 7710
rect 31164 7606 31220 7644
rect 30828 7298 30884 7308
rect 31052 7362 31108 7374
rect 31052 7310 31054 7362
rect 31106 7310 31108 7362
rect 30940 7252 30996 7262
rect 30716 6692 30772 6702
rect 30940 6692 30996 7196
rect 31052 7028 31108 7310
rect 31052 6962 31108 6972
rect 31164 7364 31220 7374
rect 30716 6690 30996 6692
rect 30716 6638 30718 6690
rect 30770 6638 30996 6690
rect 30716 6636 30996 6638
rect 30716 6626 30772 6636
rect 27804 6468 27860 6478
rect 27468 6132 27524 6142
rect 27468 6038 27524 6076
rect 27804 6130 27860 6412
rect 30380 6468 30436 6478
rect 30380 6374 30436 6412
rect 31052 6468 31108 6478
rect 31052 6374 31108 6412
rect 27804 6078 27806 6130
rect 27858 6078 27860 6130
rect 27804 6066 27860 6078
rect 27356 5854 27358 5906
rect 27410 5854 27412 5906
rect 27356 4452 27412 5854
rect 27692 5908 27748 5918
rect 27692 5814 27748 5852
rect 27580 5794 27636 5806
rect 27580 5742 27582 5794
rect 27634 5742 27636 5794
rect 27580 5460 27636 5742
rect 27580 5404 28196 5460
rect 28140 5346 28196 5404
rect 28140 5294 28142 5346
rect 28194 5294 28196 5346
rect 28140 5282 28196 5294
rect 27804 5124 27860 5134
rect 27804 5030 27860 5068
rect 28476 5124 28532 5134
rect 28476 5030 28532 5068
rect 31164 5122 31220 7308
rect 31164 5070 31166 5122
rect 31218 5070 31220 5122
rect 28252 4900 28308 4910
rect 28252 4806 28308 4844
rect 29932 4900 29988 4910
rect 27356 4396 27860 4452
rect 27804 4226 27860 4396
rect 29932 4450 29988 4844
rect 29932 4398 29934 4450
rect 29986 4398 29988 4450
rect 29932 4386 29988 4398
rect 27804 4174 27806 4226
rect 27858 4174 27860 4226
rect 27804 4162 27860 4174
rect 30604 4340 30660 4350
rect 31164 4340 31220 5070
rect 31276 5124 31332 8988
rect 31388 8978 31444 8988
rect 31612 8370 31668 9212
rect 31724 9202 31780 9212
rect 31836 9156 31892 10670
rect 33404 10388 33460 11116
rect 32172 9716 32228 9726
rect 31948 9156 32004 9166
rect 31836 9100 31948 9156
rect 31948 9062 32004 9100
rect 32172 9154 32228 9660
rect 32172 9102 32174 9154
rect 32226 9102 32228 9154
rect 32172 9090 32228 9102
rect 33068 9156 33124 9166
rect 33068 9042 33124 9100
rect 33404 9154 33460 10332
rect 33404 9102 33406 9154
rect 33458 9102 33460 9154
rect 33404 9090 33460 9102
rect 33516 10500 33572 10510
rect 33068 8990 33070 9042
rect 33122 8990 33124 9042
rect 33068 8978 33124 8990
rect 31724 8820 31780 8830
rect 31724 8726 31780 8764
rect 33068 8820 33124 8830
rect 33068 8726 33124 8764
rect 31612 8318 31614 8370
rect 31666 8318 31668 8370
rect 31612 8306 31668 8318
rect 31388 8148 31444 8158
rect 31388 6916 31444 8092
rect 31836 7700 31892 7710
rect 31836 7606 31892 7644
rect 31388 6578 31444 6860
rect 32844 6916 32900 6926
rect 32844 6822 32900 6860
rect 33516 6690 33572 10444
rect 33852 9828 33908 12124
rect 33740 9826 33908 9828
rect 33740 9774 33854 9826
rect 33906 9774 33908 9826
rect 33740 9772 33908 9774
rect 33628 9602 33684 9614
rect 33628 9550 33630 9602
rect 33682 9550 33684 9602
rect 33628 9156 33684 9550
rect 33628 9090 33684 9100
rect 33740 8370 33796 9772
rect 33852 9762 33908 9772
rect 33740 8318 33742 8370
rect 33794 8318 33796 8370
rect 33740 8306 33796 8318
rect 34188 7700 34244 16828
rect 34860 16210 34916 16222
rect 34860 16158 34862 16210
rect 34914 16158 34916 16210
rect 34300 15876 34356 15886
rect 34300 15538 34356 15820
rect 34300 15486 34302 15538
rect 34354 15486 34356 15538
rect 34300 15474 34356 15486
rect 34748 12964 34804 12974
rect 34636 12908 34748 12964
rect 34636 12850 34692 12908
rect 34748 12898 34804 12908
rect 34636 12798 34638 12850
rect 34690 12798 34692 12850
rect 34636 12786 34692 12798
rect 34300 12738 34356 12750
rect 34300 12686 34302 12738
rect 34354 12686 34356 12738
rect 34300 12404 34356 12686
rect 34860 12628 34916 16158
rect 34972 16098 35028 20524
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35420 17780 35476 17790
rect 35532 17780 35588 24668
rect 35644 23940 35700 23950
rect 35644 23846 35700 23884
rect 35980 23828 36036 23838
rect 35980 23734 36036 23772
rect 36092 23828 36148 27132
rect 36316 27076 36372 27086
rect 36316 26982 36372 27020
rect 36428 25620 36484 27692
rect 36652 26908 36708 27804
rect 36652 26852 36820 26908
rect 36428 25554 36484 25564
rect 36316 25172 36372 25182
rect 36204 24610 36260 24622
rect 36204 24558 36206 24610
rect 36258 24558 36260 24610
rect 36204 24050 36260 24558
rect 36204 23998 36206 24050
rect 36258 23998 36260 24050
rect 36204 23986 36260 23998
rect 36316 23938 36372 25116
rect 36316 23886 36318 23938
rect 36370 23886 36372 23938
rect 36316 23874 36372 23886
rect 36092 23826 36260 23828
rect 36092 23774 36094 23826
rect 36146 23774 36260 23826
rect 36092 23772 36260 23774
rect 36092 23762 36148 23772
rect 36204 23492 36260 23772
rect 36204 23436 36596 23492
rect 36540 23378 36596 23436
rect 36540 23326 36542 23378
rect 36594 23326 36596 23378
rect 36540 23314 36596 23326
rect 36764 23156 36820 26852
rect 36988 24164 37044 28252
rect 37100 27300 37156 27310
rect 37100 27206 37156 27244
rect 37212 27076 37268 27086
rect 37212 26982 37268 27020
rect 37660 26964 37716 27002
rect 37660 26898 37716 26908
rect 37100 26852 37156 26862
rect 37100 26758 37156 26796
rect 37772 26516 37828 28364
rect 37996 27524 38052 28478
rect 38108 28530 38164 28542
rect 38108 28478 38110 28530
rect 38162 28478 38164 28530
rect 38108 27748 38164 28478
rect 38108 27682 38164 27692
rect 37996 27468 38276 27524
rect 37996 26962 38052 26974
rect 37996 26910 37998 26962
rect 38050 26910 38052 26962
rect 37660 26460 37828 26516
rect 37884 26852 37940 26862
rect 36988 24108 37380 24164
rect 37212 23940 37268 23950
rect 37212 23846 37268 23884
rect 36876 23828 36932 23838
rect 36876 23734 36932 23772
rect 37100 23716 37156 23726
rect 36764 23090 36820 23100
rect 36988 23660 37100 23716
rect 36428 22146 36484 22158
rect 36428 22094 36430 22146
rect 36482 22094 36484 22146
rect 35644 21700 35700 21710
rect 35644 21476 35700 21644
rect 35644 21410 35700 21420
rect 36092 21588 36148 21598
rect 35476 17724 35588 17780
rect 35980 20692 36036 20702
rect 35980 18338 36036 20636
rect 35980 18286 35982 18338
rect 36034 18286 36036 18338
rect 35420 17714 35476 17724
rect 35980 16772 36036 18286
rect 35980 16706 36036 16716
rect 36092 16548 36148 21532
rect 36204 21476 36260 21486
rect 36204 21382 36260 21420
rect 36428 19012 36484 22094
rect 36428 18946 36484 18956
rect 36988 22148 37044 23660
rect 37100 23622 37156 23660
rect 37212 23380 37268 23390
rect 37324 23380 37380 24108
rect 37660 23604 37716 26460
rect 37772 26292 37828 26302
rect 37884 26292 37940 26796
rect 37772 26290 37940 26292
rect 37772 26238 37774 26290
rect 37826 26238 37940 26290
rect 37772 26236 37940 26238
rect 37772 26226 37828 26236
rect 37996 26066 38052 26910
rect 37996 26014 37998 26066
rect 38050 26014 38052 26066
rect 37996 24836 38052 26014
rect 37996 24770 38052 24780
rect 37996 24612 38052 24622
rect 37660 23548 37940 23604
rect 37772 23380 37828 23390
rect 37212 23378 37828 23380
rect 37212 23326 37214 23378
rect 37266 23326 37774 23378
rect 37826 23326 37828 23378
rect 37212 23324 37828 23326
rect 37212 23314 37268 23324
rect 37100 23154 37156 23166
rect 37100 23102 37102 23154
rect 37154 23102 37156 23154
rect 37100 22484 37156 23102
rect 37212 22932 37268 22942
rect 37212 22838 37268 22876
rect 37100 22418 37156 22428
rect 37324 22258 37380 22270
rect 37324 22206 37326 22258
rect 37378 22206 37380 22258
rect 37324 22148 37380 22206
rect 36988 22092 37380 22148
rect 36988 18452 37044 22092
rect 37436 22036 37492 23324
rect 37772 23314 37828 23324
rect 37212 21980 37492 22036
rect 37100 21586 37156 21598
rect 37100 21534 37102 21586
rect 37154 21534 37156 21586
rect 37100 21364 37156 21534
rect 37100 21298 37156 21308
rect 37212 20132 37268 21980
rect 37772 21588 37828 21598
rect 37772 20916 37828 21532
rect 37772 20850 37828 20860
rect 37660 20804 37716 20814
rect 37548 20748 37660 20804
rect 37324 20692 37380 20702
rect 37324 20598 37380 20636
rect 37436 20132 37492 20142
rect 37548 20132 37604 20748
rect 37660 20738 37716 20748
rect 37884 20132 37940 23548
rect 37996 22370 38052 24556
rect 37996 22318 37998 22370
rect 38050 22318 38052 22370
rect 37996 20802 38052 22318
rect 38108 23492 38164 23502
rect 38108 21586 38164 23436
rect 38108 21534 38110 21586
rect 38162 21534 38164 21586
rect 38108 21522 38164 21534
rect 37996 20750 37998 20802
rect 38050 20750 38052 20802
rect 37996 20738 38052 20750
rect 37212 20130 37380 20132
rect 37212 20078 37214 20130
rect 37266 20078 37380 20130
rect 37212 20076 37380 20078
rect 37212 20066 37268 20076
rect 37100 20018 37156 20030
rect 37100 19966 37102 20018
rect 37154 19966 37156 20018
rect 37100 19908 37156 19966
rect 37100 19842 37156 19852
rect 37324 19796 37380 20076
rect 37436 20130 37604 20132
rect 37436 20078 37438 20130
rect 37490 20078 37604 20130
rect 37436 20076 37604 20078
rect 37772 20076 37940 20132
rect 37436 20066 37492 20076
rect 37548 19796 37604 19806
rect 37324 19794 37604 19796
rect 37324 19742 37550 19794
rect 37602 19742 37604 19794
rect 37324 19740 37604 19742
rect 37548 19730 37604 19740
rect 37772 19460 37828 20076
rect 37884 19906 37940 19918
rect 37884 19854 37886 19906
rect 37938 19854 37940 19906
rect 37884 19794 37940 19854
rect 37884 19742 37886 19794
rect 37938 19742 37940 19794
rect 37884 19730 37940 19742
rect 37772 19394 37828 19404
rect 37212 19346 37268 19358
rect 38220 19348 38276 27468
rect 38332 26292 38388 32508
rect 38444 31890 38500 33628
rect 38668 32788 38724 32798
rect 38668 32694 38724 32732
rect 38780 32340 38836 34300
rect 38892 34916 38948 34926
rect 39116 34916 39172 34926
rect 38892 34914 39116 34916
rect 38892 34862 38894 34914
rect 38946 34862 39116 34914
rect 38892 34860 39116 34862
rect 38892 34130 38948 34860
rect 39116 34850 39172 34860
rect 39228 34914 39284 34972
rect 39228 34862 39230 34914
rect 39282 34862 39284 34914
rect 39228 34850 39284 34862
rect 39004 34692 39060 34702
rect 39004 34598 39060 34636
rect 39116 34692 39172 34702
rect 39340 34692 39396 35644
rect 39452 35634 39508 35644
rect 39788 35588 39844 35598
rect 39676 35586 39844 35588
rect 39676 35534 39790 35586
rect 39842 35534 39844 35586
rect 39676 35532 39844 35534
rect 39676 35308 39732 35532
rect 39788 35522 39844 35532
rect 39116 34690 39396 34692
rect 39116 34638 39118 34690
rect 39170 34638 39396 34690
rect 39116 34636 39396 34638
rect 39452 35252 39732 35308
rect 39452 34802 39508 35252
rect 39788 34916 39844 34926
rect 40012 34916 40068 38612
rect 40236 36932 40292 38894
rect 40460 38836 40516 38846
rect 40796 38836 40852 38846
rect 40460 38834 40852 38836
rect 40460 38782 40462 38834
rect 40514 38782 40798 38834
rect 40850 38782 40852 38834
rect 40460 38780 40852 38782
rect 40460 38770 40516 38780
rect 40796 38770 40852 38780
rect 41132 38668 41188 39006
rect 41244 38946 41300 39228
rect 41244 38894 41246 38946
rect 41298 38894 41300 38946
rect 41244 38882 41300 38894
rect 41356 38836 41412 38846
rect 41356 38742 41412 38780
rect 41132 38612 41412 38668
rect 41356 38162 41412 38612
rect 41356 38110 41358 38162
rect 41410 38110 41412 38162
rect 41356 38098 41412 38110
rect 40236 36820 40292 36876
rect 40236 36764 40740 36820
rect 40572 36484 40628 36494
rect 40572 36390 40628 36428
rect 40684 36370 40740 36764
rect 40684 36318 40686 36370
rect 40738 36318 40740 36370
rect 40684 36306 40740 36318
rect 40908 36260 40964 36270
rect 40908 36258 41748 36260
rect 40908 36206 40910 36258
rect 40962 36206 41748 36258
rect 40908 36204 41748 36206
rect 40908 36194 40964 36204
rect 40236 35924 40292 35934
rect 40124 35364 40180 35374
rect 40124 35026 40180 35308
rect 40124 34974 40126 35026
rect 40178 34974 40180 35026
rect 40124 34962 40180 34974
rect 39844 34860 39956 34916
rect 39788 34822 39844 34860
rect 39452 34750 39454 34802
rect 39506 34750 39508 34802
rect 39116 34626 39172 34636
rect 38892 34078 38894 34130
rect 38946 34078 38948 34130
rect 38892 32562 38948 34078
rect 39228 32900 39284 32910
rect 39116 32788 39172 32798
rect 39116 32694 39172 32732
rect 39228 32786 39284 32844
rect 39228 32734 39230 32786
rect 39282 32734 39284 32786
rect 39228 32722 39284 32734
rect 38892 32510 38894 32562
rect 38946 32510 38948 32562
rect 38892 32498 38948 32510
rect 39340 32562 39396 32574
rect 39340 32510 39342 32562
rect 39394 32510 39396 32562
rect 39340 32452 39396 32510
rect 38780 32284 38948 32340
rect 38444 31838 38446 31890
rect 38498 31838 38500 31890
rect 38444 31826 38500 31838
rect 38780 29314 38836 29326
rect 38780 29262 38782 29314
rect 38834 29262 38836 29314
rect 38780 28644 38836 29262
rect 38780 28578 38836 28588
rect 38892 28084 38948 32284
rect 39228 32004 39284 32014
rect 39004 31948 39228 32004
rect 39004 31778 39060 31948
rect 39004 31726 39006 31778
rect 39058 31726 39060 31778
rect 39004 31714 39060 31726
rect 39004 30884 39060 30894
rect 39004 28644 39060 30828
rect 39116 29428 39172 31948
rect 39228 31938 39284 31948
rect 39228 31780 39284 31790
rect 39228 29652 39284 31724
rect 39340 29764 39396 32396
rect 39452 30212 39508 34750
rect 39564 34468 39620 34478
rect 39564 34354 39620 34412
rect 39564 34302 39566 34354
rect 39618 34302 39620 34354
rect 39564 34290 39620 34302
rect 39900 33348 39956 34860
rect 40012 34850 40068 34860
rect 40236 34916 40292 35868
rect 40908 35810 40964 35822
rect 40908 35758 40910 35810
rect 40962 35758 40964 35810
rect 40236 34850 40292 34860
rect 40348 35588 40404 35598
rect 40908 35588 40964 35758
rect 41244 35812 41300 35822
rect 41132 35700 41188 35710
rect 41244 35700 41300 35756
rect 41132 35698 41300 35700
rect 41132 35646 41134 35698
rect 41186 35646 41300 35698
rect 41132 35644 41300 35646
rect 41132 35634 41188 35644
rect 40348 35586 40964 35588
rect 40348 35534 40350 35586
rect 40402 35534 40964 35586
rect 40348 35532 40964 35534
rect 40012 34690 40068 34702
rect 40012 34638 40014 34690
rect 40066 34638 40068 34690
rect 40012 34468 40068 34638
rect 40236 34692 40292 34702
rect 40236 34598 40292 34636
rect 40012 34402 40068 34412
rect 39900 33292 40068 33348
rect 39900 33122 39956 33134
rect 39900 33070 39902 33122
rect 39954 33070 39956 33122
rect 39900 33012 39956 33070
rect 39788 32956 39956 33012
rect 39564 32564 39620 32574
rect 39788 32564 39844 32956
rect 39900 32788 39956 32798
rect 40012 32788 40068 33292
rect 39900 32786 40068 32788
rect 39900 32734 39902 32786
rect 39954 32734 40068 32786
rect 39900 32732 40068 32734
rect 39900 32722 39956 32732
rect 39564 32562 39844 32564
rect 39564 32510 39566 32562
rect 39618 32510 39844 32562
rect 39564 32508 39844 32510
rect 40124 32562 40180 32574
rect 40124 32510 40126 32562
rect 40178 32510 40180 32562
rect 39564 31556 39620 32508
rect 40124 32004 40180 32510
rect 40124 31938 40180 31948
rect 39900 31780 39956 31790
rect 39900 31686 39956 31724
rect 39564 31490 39620 31500
rect 40348 31220 40404 35532
rect 40460 34802 40516 34814
rect 40460 34750 40462 34802
rect 40514 34750 40516 34802
rect 40460 34692 40516 34750
rect 41020 34692 41076 34702
rect 40460 34690 41076 34692
rect 40460 34638 41022 34690
rect 41074 34638 41076 34690
rect 40460 34636 41076 34638
rect 40460 31444 40516 34636
rect 41020 34626 41076 34636
rect 41244 33124 41300 35644
rect 41692 35698 41748 36204
rect 41692 35646 41694 35698
rect 41746 35646 41748 35698
rect 41692 35634 41748 35646
rect 41580 34914 41636 34926
rect 41580 34862 41582 34914
rect 41634 34862 41636 34914
rect 41580 34804 41636 34862
rect 41580 34738 41636 34748
rect 41244 33058 41300 33068
rect 41580 34020 41636 34030
rect 41580 33012 41636 33964
rect 41692 33348 41748 33358
rect 41692 33254 41748 33292
rect 41580 32946 41636 32956
rect 41804 32788 41860 43652
rect 41916 43426 41972 45052
rect 42476 45108 42532 45166
rect 42476 45042 42532 45052
rect 42364 44994 42420 45006
rect 42364 44942 42366 44994
rect 42418 44942 42420 44994
rect 42140 44436 42196 44446
rect 42364 44436 42420 44942
rect 42140 44434 42420 44436
rect 42140 44382 42142 44434
rect 42194 44382 42420 44434
rect 42140 44380 42420 44382
rect 42140 44370 42196 44380
rect 42588 43540 42644 45612
rect 44268 45666 44324 45678
rect 44268 45614 44270 45666
rect 44322 45614 44324 45666
rect 43820 45332 43876 45342
rect 43708 45220 43764 45230
rect 43820 45220 43876 45276
rect 44268 45332 44324 45614
rect 44268 45266 44324 45276
rect 43708 45218 43876 45220
rect 43708 45166 43710 45218
rect 43762 45166 43876 45218
rect 43708 45164 43876 45166
rect 44156 45220 44212 45230
rect 43708 44996 43764 45164
rect 43708 44930 43764 44940
rect 44156 44436 44212 45164
rect 45276 44994 45332 46620
rect 45276 44942 45278 44994
rect 45330 44942 45332 44994
rect 45276 44930 45332 44942
rect 45388 46002 45444 46014
rect 45388 45950 45390 46002
rect 45442 45950 45444 46002
rect 44268 44436 44324 44446
rect 44156 44434 44324 44436
rect 44156 44382 44270 44434
rect 44322 44382 44324 44434
rect 44156 44380 44324 44382
rect 44268 44212 44324 44380
rect 45052 44324 45108 44334
rect 45052 44230 45108 44268
rect 44268 44146 44324 44156
rect 44940 44212 44996 44222
rect 44940 44118 44996 44156
rect 44716 44098 44772 44110
rect 44716 44046 44718 44098
rect 44770 44046 44772 44098
rect 43708 43764 43764 43774
rect 42588 43474 42644 43484
rect 43484 43652 43540 43662
rect 41916 43374 41918 43426
rect 41970 43374 41972 43426
rect 41916 42308 41972 43374
rect 41916 42242 41972 42252
rect 42588 41300 42644 41310
rect 41916 40516 41972 40526
rect 41916 40180 41972 40460
rect 42028 40404 42084 40414
rect 42028 40310 42084 40348
rect 41916 40124 42084 40180
rect 42028 37492 42084 40124
rect 42140 38052 42196 38062
rect 42588 38052 42644 41244
rect 43036 41298 43092 41310
rect 43036 41246 43038 41298
rect 43090 41246 43092 41298
rect 43036 40516 43092 41246
rect 43484 41300 43540 43596
rect 43484 41206 43540 41244
rect 43036 40450 43092 40460
rect 43148 40964 43204 40974
rect 42140 38050 42644 38052
rect 42140 37998 42142 38050
rect 42194 37998 42644 38050
rect 42140 37996 42644 37998
rect 42140 37986 42196 37996
rect 42588 37826 42644 37996
rect 42588 37774 42590 37826
rect 42642 37774 42644 37826
rect 42028 37436 42308 37492
rect 42252 36370 42308 37436
rect 42588 37268 42644 37774
rect 42924 37268 42980 37278
rect 42588 37266 42980 37268
rect 42588 37214 42926 37266
rect 42978 37214 42980 37266
rect 42588 37212 42980 37214
rect 42924 37202 42980 37212
rect 43036 36484 43092 36494
rect 42252 36318 42254 36370
rect 42306 36318 42308 36370
rect 42252 36306 42308 36318
rect 42364 36370 42420 36382
rect 42364 36318 42366 36370
rect 42418 36318 42420 36370
rect 42028 36258 42084 36270
rect 42028 36206 42030 36258
rect 42082 36206 42084 36258
rect 42028 34356 42084 36206
rect 42364 35812 42420 36318
rect 42252 35756 42420 35812
rect 42924 36258 42980 36270
rect 42924 36206 42926 36258
rect 42978 36206 42980 36258
rect 42924 35812 42980 36206
rect 43036 35922 43092 36428
rect 43036 35870 43038 35922
rect 43090 35870 43092 35922
rect 43036 35858 43092 35870
rect 42140 35700 42196 35710
rect 42140 35606 42196 35644
rect 42252 34804 42308 35756
rect 42924 35746 42980 35756
rect 42700 35700 42756 35710
rect 42252 34738 42308 34748
rect 42364 35698 42756 35700
rect 42364 35646 42702 35698
rect 42754 35646 42756 35698
rect 42364 35644 42756 35646
rect 42140 34690 42196 34702
rect 42140 34638 42142 34690
rect 42194 34638 42196 34690
rect 42140 34468 42196 34638
rect 42364 34468 42420 35644
rect 42700 35634 42756 35644
rect 42476 35476 42532 35486
rect 42812 35476 42868 35486
rect 42476 35474 42812 35476
rect 42476 35422 42478 35474
rect 42530 35422 42812 35474
rect 42476 35420 42812 35422
rect 42476 35410 42532 35420
rect 42812 35410 42868 35420
rect 43148 35252 43204 40908
rect 43708 40404 43764 43708
rect 44716 43708 44772 44046
rect 45276 44098 45332 44110
rect 45276 44046 45278 44098
rect 45330 44046 45332 44098
rect 44492 43652 44548 43662
rect 44716 43652 44884 43708
rect 44492 43558 44548 43596
rect 44604 41858 44660 41870
rect 44604 41806 44606 41858
rect 44658 41806 44660 41858
rect 44604 41412 44660 41806
rect 44268 41356 44660 41412
rect 44044 41074 44100 41086
rect 44044 41022 44046 41074
rect 44098 41022 44100 41074
rect 43596 40348 43764 40404
rect 43932 40516 43988 40526
rect 43596 35476 43652 40348
rect 43708 39060 43764 39070
rect 43708 37378 43764 39004
rect 43708 37326 43710 37378
rect 43762 37326 43764 37378
rect 43708 37314 43764 37326
rect 43820 38836 43876 38846
rect 43708 36484 43764 36494
rect 43708 36390 43764 36428
rect 43820 36370 43876 38780
rect 43932 37940 43988 40460
rect 44044 40404 44100 41022
rect 44156 40964 44212 40974
rect 44268 40964 44324 41356
rect 44380 41188 44436 41198
rect 44716 41188 44772 41198
rect 44380 41186 44772 41188
rect 44380 41134 44382 41186
rect 44434 41134 44718 41186
rect 44770 41134 44772 41186
rect 44380 41132 44772 41134
rect 44380 41122 44436 41132
rect 44716 41122 44772 41132
rect 44212 40908 44324 40964
rect 44156 40870 44212 40908
rect 44044 39508 44100 40348
rect 44828 39732 44884 43652
rect 44940 42084 44996 42094
rect 44940 40740 44996 42028
rect 45052 41860 45108 41870
rect 45052 40962 45108 41804
rect 45164 41188 45220 41198
rect 45276 41188 45332 44046
rect 45388 43652 45444 45950
rect 45500 44210 45556 47404
rect 45836 49026 46116 49028
rect 45836 48974 46062 49026
rect 46114 48974 46116 49026
rect 45836 48972 46116 48974
rect 45836 46340 45892 48972
rect 46060 48962 46116 48972
rect 45948 48804 46004 48814
rect 46396 48804 46452 48814
rect 45948 48802 46452 48804
rect 45948 48750 45950 48802
rect 46002 48750 46398 48802
rect 46450 48750 46452 48802
rect 45948 48748 46452 48750
rect 45948 48738 46004 48748
rect 46284 48242 46340 48254
rect 46284 48190 46286 48242
rect 46338 48190 46340 48242
rect 45948 48132 46004 48142
rect 46284 48132 46340 48190
rect 45948 48130 46340 48132
rect 45948 48078 45950 48130
rect 46002 48078 46340 48130
rect 45948 48076 46340 48078
rect 46396 48132 46452 48748
rect 46508 48468 46564 50430
rect 48636 49028 48692 50654
rect 49196 50596 49252 50606
rect 49084 50540 49196 50596
rect 48748 49980 49028 50036
rect 48748 49250 48804 49980
rect 48972 49924 49028 49980
rect 48972 49830 49028 49868
rect 48860 49812 48916 49822
rect 48860 49718 48916 49756
rect 48972 49588 49028 49598
rect 49084 49588 49140 50540
rect 49196 50530 49252 50540
rect 49756 50596 49812 50606
rect 49196 50370 49252 50382
rect 49196 50318 49198 50370
rect 49250 50318 49252 50370
rect 49196 49812 49252 50318
rect 49756 50034 49812 50540
rect 49756 49982 49758 50034
rect 49810 49982 49812 50034
rect 49756 49970 49812 49982
rect 49868 50034 49924 51324
rect 51100 50818 51156 51548
rect 51100 50766 51102 50818
rect 51154 50766 51156 50818
rect 51100 50754 51156 50766
rect 51212 51378 51268 51390
rect 51212 51326 51214 51378
rect 51266 51326 51268 51378
rect 49868 49982 49870 50034
rect 49922 49982 49924 50034
rect 49868 49970 49924 49982
rect 49980 50484 50036 50494
rect 49980 50034 50036 50428
rect 51212 50484 51268 51326
rect 51436 51378 51492 51390
rect 51436 51326 51438 51378
rect 51490 51326 51492 51378
rect 51212 50418 51268 50428
rect 51324 51266 51380 51278
rect 51324 51214 51326 51266
rect 51378 51214 51380 51266
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 49980 49982 49982 50034
rect 50034 49982 50036 50034
rect 49420 49812 49476 49822
rect 49196 49810 49476 49812
rect 49196 49758 49422 49810
rect 49474 49758 49476 49810
rect 49196 49756 49476 49758
rect 48972 49586 49140 49588
rect 48972 49534 48974 49586
rect 49026 49534 49140 49586
rect 48972 49532 49140 49534
rect 48972 49522 49028 49532
rect 48748 49198 48750 49250
rect 48802 49198 48804 49250
rect 48748 49186 48804 49198
rect 48972 49028 49028 49038
rect 49196 49028 49252 49038
rect 48636 49026 49028 49028
rect 48636 48974 48974 49026
rect 49026 48974 49028 49026
rect 48636 48972 49028 48974
rect 46620 48804 46676 48814
rect 46620 48710 46676 48748
rect 46732 48802 46788 48814
rect 46732 48750 46734 48802
rect 46786 48750 46788 48802
rect 46620 48468 46676 48478
rect 46508 48466 46676 48468
rect 46508 48414 46622 48466
rect 46674 48414 46676 48466
rect 46508 48412 46676 48414
rect 46620 48402 46676 48412
rect 46732 48356 46788 48750
rect 47180 48804 47236 48814
rect 46844 48356 46900 48366
rect 46732 48354 46900 48356
rect 46732 48302 46846 48354
rect 46898 48302 46900 48354
rect 46732 48300 46900 48302
rect 46844 48290 46900 48300
rect 47180 48356 47236 48748
rect 47180 48262 47236 48300
rect 48300 48802 48356 48814
rect 48300 48750 48302 48802
rect 48354 48750 48356 48802
rect 46620 48242 46676 48254
rect 46620 48190 46622 48242
rect 46674 48190 46676 48242
rect 46508 48132 46564 48142
rect 46396 48076 46508 48132
rect 45948 47124 46004 48076
rect 46508 48066 46564 48076
rect 46620 48020 46676 48190
rect 46620 47954 46676 47964
rect 47404 48132 47460 48142
rect 47404 48018 47460 48076
rect 48188 48132 48244 48142
rect 48188 48038 48244 48076
rect 47404 47966 47406 48018
rect 47458 47966 47460 48018
rect 46844 47234 46900 47246
rect 46844 47182 46846 47234
rect 46898 47182 46900 47234
rect 46844 47124 46900 47182
rect 47404 47124 47460 47966
rect 47740 48020 47796 48030
rect 47740 47460 47796 47964
rect 47740 47394 47796 47404
rect 46844 47068 47460 47124
rect 45948 47058 46004 47068
rect 45836 46274 45892 46284
rect 46284 46562 46340 46574
rect 46284 46510 46286 46562
rect 46338 46510 46340 46562
rect 46284 45668 46340 46510
rect 46060 45612 46284 45668
rect 45612 44324 45668 44334
rect 45948 44324 46004 44334
rect 45668 44322 46004 44324
rect 45668 44270 45950 44322
rect 46002 44270 46004 44322
rect 45668 44268 46004 44270
rect 45612 44230 45668 44268
rect 45948 44258 46004 44268
rect 45500 44158 45502 44210
rect 45554 44158 45556 44210
rect 45500 44146 45556 44158
rect 46060 44210 46116 45612
rect 46284 45602 46340 45612
rect 47068 45890 47124 45902
rect 47068 45838 47070 45890
rect 47122 45838 47124 45890
rect 46620 45332 46676 45342
rect 47068 45332 47124 45838
rect 46676 45276 47124 45332
rect 46620 45106 46676 45276
rect 46620 45054 46622 45106
rect 46674 45054 46676 45106
rect 46620 45042 46676 45054
rect 47068 44884 47124 44894
rect 47180 44884 47236 47068
rect 47852 46786 47908 46798
rect 47852 46734 47854 46786
rect 47906 46734 47908 46786
rect 47740 46674 47796 46686
rect 47740 46622 47742 46674
rect 47794 46622 47796 46674
rect 47740 46340 47796 46622
rect 47740 46274 47796 46284
rect 47740 45780 47796 45790
rect 47124 44828 47236 44884
rect 47292 45778 47796 45780
rect 47292 45726 47742 45778
rect 47794 45726 47796 45778
rect 47292 45724 47796 45726
rect 47068 44818 47124 44828
rect 46060 44158 46062 44210
rect 46114 44158 46116 44210
rect 46060 44146 46116 44158
rect 46284 44098 46340 44110
rect 46284 44046 46286 44098
rect 46338 44046 46340 44098
rect 45388 43586 45444 43596
rect 46060 43652 46116 43662
rect 45164 41186 45332 41188
rect 45164 41134 45166 41186
rect 45218 41134 45332 41186
rect 45164 41132 45332 41134
rect 45164 41122 45220 41132
rect 45388 41076 45444 41086
rect 45388 41074 45556 41076
rect 45388 41022 45390 41074
rect 45442 41022 45556 41074
rect 45388 41020 45556 41022
rect 45388 41010 45444 41020
rect 45052 40910 45054 40962
rect 45106 40910 45108 40962
rect 45052 40898 45108 40910
rect 44940 40684 45332 40740
rect 44940 40402 44996 40414
rect 44940 40350 44942 40402
rect 44994 40350 44996 40402
rect 44940 39842 44996 40350
rect 45276 40402 45332 40684
rect 45276 40350 45278 40402
rect 45330 40350 45332 40402
rect 45276 40338 45332 40350
rect 45500 40402 45556 41020
rect 45500 40350 45502 40402
rect 45554 40350 45556 40402
rect 45164 40292 45220 40302
rect 45164 40198 45220 40236
rect 44940 39790 44942 39842
rect 44994 39790 44996 39842
rect 44940 39778 44996 39790
rect 44044 39442 44100 39452
rect 44492 39676 44884 39732
rect 44380 39060 44436 39098
rect 44380 38994 44436 39004
rect 44044 38834 44100 38846
rect 44044 38782 44046 38834
rect 44098 38782 44100 38834
rect 44044 38724 44100 38782
rect 44380 38836 44436 38846
rect 44492 38836 44548 39676
rect 44828 39508 44884 39518
rect 44828 38948 44884 39452
rect 44940 39394 44996 39406
rect 44940 39342 44942 39394
rect 44994 39342 44996 39394
rect 44940 39172 44996 39342
rect 44940 39106 44996 39116
rect 44940 38948 44996 38958
rect 44828 38946 44996 38948
rect 44828 38894 44942 38946
rect 44994 38894 44996 38946
rect 44828 38892 44996 38894
rect 44940 38882 44996 38892
rect 45052 38948 45108 38958
rect 45052 38946 45220 38948
rect 45052 38894 45054 38946
rect 45106 38894 45220 38946
rect 45052 38892 45220 38894
rect 45052 38882 45108 38892
rect 44380 38834 44548 38836
rect 44380 38782 44382 38834
rect 44434 38782 44548 38834
rect 44380 38780 44548 38782
rect 44716 38836 44772 38846
rect 44716 38834 44884 38836
rect 44716 38782 44718 38834
rect 44770 38782 44884 38834
rect 44716 38780 44884 38782
rect 44380 38770 44436 38780
rect 44716 38770 44772 38780
rect 44044 38658 44100 38668
rect 44828 38668 44884 38780
rect 44828 38612 45108 38668
rect 45052 38610 45108 38612
rect 45052 38558 45054 38610
rect 45106 38558 45108 38610
rect 45052 38546 45108 38558
rect 43932 37884 44548 37940
rect 43820 36318 43822 36370
rect 43874 36318 43876 36370
rect 43820 36306 43876 36318
rect 44380 37716 44436 37726
rect 44044 36258 44100 36270
rect 44268 36260 44324 36270
rect 44044 36206 44046 36258
rect 44098 36206 44100 36258
rect 43596 35410 43652 35420
rect 43708 35698 43764 35710
rect 43708 35646 43710 35698
rect 43762 35646 43764 35698
rect 43708 35364 43764 35646
rect 43708 35298 43764 35308
rect 43932 35698 43988 35710
rect 43932 35646 43934 35698
rect 43986 35646 43988 35698
rect 43932 35364 43988 35646
rect 43932 35298 43988 35308
rect 42588 35196 43204 35252
rect 43372 35252 43428 35262
rect 42476 34804 42532 34814
rect 42476 34710 42532 34748
rect 42588 34802 42644 35196
rect 42588 34750 42590 34802
rect 42642 34750 42644 34802
rect 42588 34738 42644 34750
rect 42812 34692 42868 34702
rect 42140 34412 42420 34468
rect 42028 34300 42308 34356
rect 42028 33348 42084 33358
rect 42028 33234 42084 33292
rect 42028 33182 42030 33234
rect 42082 33182 42084 33234
rect 42028 33170 42084 33182
rect 42140 33346 42196 33358
rect 42140 33294 42142 33346
rect 42194 33294 42196 33346
rect 42140 33124 42196 33294
rect 42140 33058 42196 33068
rect 41244 32732 41860 32788
rect 42252 32786 42308 34300
rect 42252 32734 42254 32786
rect 42306 32734 42308 32786
rect 40572 31668 40628 31678
rect 40572 31666 41188 31668
rect 40572 31614 40574 31666
rect 40626 31614 41188 31666
rect 40572 31612 41188 31614
rect 40572 31602 40628 31612
rect 40460 31388 40964 31444
rect 40348 31154 40404 31164
rect 39452 30156 39620 30212
rect 39452 29988 39508 29998
rect 39452 29894 39508 29932
rect 39340 29698 39396 29708
rect 39228 29558 39284 29596
rect 39116 29372 39284 29428
rect 39004 28578 39060 28588
rect 39004 28418 39060 28430
rect 39004 28366 39006 28418
rect 39058 28366 39060 28418
rect 39004 28308 39060 28366
rect 39004 28242 39060 28252
rect 39116 28084 39172 28094
rect 38892 28028 39116 28084
rect 39116 28018 39172 28028
rect 38556 27748 38612 27758
rect 38444 27074 38500 27086
rect 38444 27022 38446 27074
rect 38498 27022 38500 27074
rect 38444 26964 38500 27022
rect 38444 26898 38500 26908
rect 38556 26964 38612 27692
rect 39116 27074 39172 27086
rect 39116 27022 39118 27074
rect 39170 27022 39172 27074
rect 38668 26964 38724 26974
rect 38556 26962 38724 26964
rect 38556 26910 38670 26962
rect 38722 26910 38724 26962
rect 38556 26908 38724 26910
rect 38332 26236 38500 26292
rect 38332 26068 38388 26078
rect 38332 25620 38388 26012
rect 38332 25554 38388 25564
rect 38332 24610 38388 24622
rect 38332 24558 38334 24610
rect 38386 24558 38388 24610
rect 38332 23716 38388 24558
rect 38332 23650 38388 23660
rect 38444 23492 38500 26236
rect 38556 23940 38612 26908
rect 38668 26898 38724 26908
rect 39116 26964 39172 27022
rect 39116 26898 39172 26908
rect 39228 27076 39284 29372
rect 39340 28530 39396 28542
rect 39340 28478 39342 28530
rect 39394 28478 39396 28530
rect 39340 27748 39396 28478
rect 39452 28420 39508 28430
rect 39564 28420 39620 30156
rect 40572 29988 40628 29998
rect 40348 29932 40572 29988
rect 40124 29540 40180 29550
rect 40124 29538 40292 29540
rect 40124 29486 40126 29538
rect 40178 29486 40292 29538
rect 40124 29484 40292 29486
rect 40124 29474 40180 29484
rect 39676 29426 39732 29438
rect 39676 29374 39678 29426
rect 39730 29374 39732 29426
rect 39676 28642 39732 29374
rect 39900 29316 39956 29326
rect 39900 29222 39956 29260
rect 39676 28590 39678 28642
rect 39730 28590 39732 28642
rect 39676 28578 39732 28590
rect 40012 29092 40068 29102
rect 39452 28418 39620 28420
rect 39452 28366 39454 28418
rect 39506 28366 39620 28418
rect 39452 28364 39620 28366
rect 39452 28308 39508 28364
rect 39452 28242 39508 28252
rect 39340 27682 39396 27692
rect 39564 28084 39620 28094
rect 38780 24724 38836 24734
rect 38780 24050 38836 24668
rect 39004 24724 39060 24734
rect 39004 24630 39060 24668
rect 38780 23998 38782 24050
rect 38834 23998 38836 24050
rect 38780 23986 38836 23998
rect 38556 23874 38612 23884
rect 38444 23436 38836 23492
rect 38668 21812 38724 21822
rect 38668 21586 38724 21756
rect 38668 21534 38670 21586
rect 38722 21534 38724 21586
rect 38668 21522 38724 21534
rect 37212 19294 37214 19346
rect 37266 19294 37268 19346
rect 37100 18452 37156 18462
rect 36988 18450 37156 18452
rect 36988 18398 37102 18450
rect 37154 18398 37156 18450
rect 36988 18396 37156 18398
rect 37100 18386 37156 18396
rect 36540 17780 36596 17790
rect 36540 17686 36596 17724
rect 36428 17444 36484 17454
rect 36428 17106 36484 17388
rect 36652 17220 36708 17230
rect 36428 17054 36430 17106
rect 36482 17054 36484 17106
rect 36428 17042 36484 17054
rect 36540 17164 36652 17220
rect 36316 16882 36372 16894
rect 36316 16830 36318 16882
rect 36370 16830 36372 16882
rect 36316 16772 36372 16830
rect 36316 16706 36372 16716
rect 35196 16492 35460 16502
rect 36092 16492 36372 16548
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34972 16046 34974 16098
rect 35026 16046 35028 16098
rect 34972 16034 35028 16046
rect 35644 15986 35700 15998
rect 35644 15934 35646 15986
rect 35698 15934 35700 15986
rect 35308 15540 35364 15550
rect 35308 15446 35364 15484
rect 35644 15316 35700 15934
rect 36204 15876 36260 15886
rect 35644 15250 35700 15260
rect 36092 15314 36148 15326
rect 36092 15262 36094 15314
rect 36146 15262 36148 15314
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 36092 14754 36148 15262
rect 36092 14702 36094 14754
rect 36146 14702 36148 14754
rect 35980 14418 36036 14430
rect 35980 14366 35982 14418
rect 36034 14366 36036 14418
rect 35980 13860 36036 14366
rect 35532 13804 35980 13860
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35420 13076 35476 13086
rect 35532 13076 35588 13804
rect 35980 13794 36036 13804
rect 36092 13746 36148 14702
rect 36092 13694 36094 13746
rect 36146 13694 36148 13746
rect 36092 13682 36148 13694
rect 35756 13634 35812 13646
rect 35756 13582 35758 13634
rect 35810 13582 35812 13634
rect 35420 13074 35588 13076
rect 35420 13022 35422 13074
rect 35474 13022 35588 13074
rect 35420 13020 35588 13022
rect 35644 13076 35700 13086
rect 35756 13076 35812 13582
rect 35756 13020 35924 13076
rect 35420 13010 35476 13020
rect 35644 12964 35700 13020
rect 35644 12908 35812 12964
rect 35532 12852 35588 12862
rect 34860 12562 34916 12572
rect 35308 12850 35700 12852
rect 35308 12798 35534 12850
rect 35586 12798 35700 12850
rect 35308 12796 35700 12798
rect 35084 12404 35140 12414
rect 34300 12402 35140 12404
rect 34300 12350 35086 12402
rect 35138 12350 35140 12402
rect 34300 12348 35140 12350
rect 34300 11396 34356 12348
rect 35084 12338 35140 12348
rect 35308 12402 35364 12796
rect 35532 12786 35588 12796
rect 35644 12740 35700 12796
rect 35756 12850 35812 12908
rect 35756 12798 35758 12850
rect 35810 12798 35812 12850
rect 35756 12786 35812 12798
rect 35644 12674 35700 12684
rect 35308 12350 35310 12402
rect 35362 12350 35364 12402
rect 35308 12338 35364 12350
rect 35420 12404 35476 12414
rect 35868 12404 35924 13020
rect 35420 12402 35924 12404
rect 35420 12350 35422 12402
rect 35474 12350 35924 12402
rect 35420 12348 35924 12350
rect 35420 12338 35476 12348
rect 34748 12180 34804 12190
rect 34748 12086 34804 12124
rect 35868 12178 35924 12348
rect 35980 12962 36036 12974
rect 35980 12910 35982 12962
rect 36034 12910 36036 12962
rect 35980 12404 36036 12910
rect 35980 12338 36036 12348
rect 36092 12852 36148 12862
rect 36092 12402 36148 12796
rect 36092 12350 36094 12402
rect 36146 12350 36148 12402
rect 36092 12338 36148 12350
rect 36204 12740 36260 15820
rect 36204 12402 36260 12684
rect 36316 12516 36372 16492
rect 36428 15540 36484 15550
rect 36428 15428 36484 15484
rect 36540 15428 36596 17164
rect 36652 17154 36708 17164
rect 36428 15426 36596 15428
rect 36428 15374 36430 15426
rect 36482 15374 36596 15426
rect 36428 15372 36596 15374
rect 36428 15362 36484 15372
rect 36652 13748 36708 13758
rect 36652 13654 36708 13692
rect 36428 12740 36484 12750
rect 36428 12646 36484 12684
rect 36316 12460 36484 12516
rect 36204 12350 36206 12402
rect 36258 12350 36260 12402
rect 36204 12338 36260 12350
rect 36316 12292 36372 12302
rect 36316 12198 36372 12236
rect 35868 12126 35870 12178
rect 35922 12126 35924 12178
rect 35868 12114 35924 12126
rect 35980 12178 36036 12190
rect 35980 12126 35982 12178
rect 36034 12126 36036 12178
rect 35196 12068 35252 12078
rect 34300 11330 34356 11340
rect 35084 12012 35196 12068
rect 35084 11284 35140 12012
rect 35196 12002 35252 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 9044 35140 11228
rect 35644 10948 35700 10958
rect 35644 10610 35700 10892
rect 35868 10836 35924 10846
rect 35644 10558 35646 10610
rect 35698 10558 35700 10610
rect 35644 10546 35700 10558
rect 35756 10724 35812 10734
rect 35644 10388 35700 10398
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 9604 35588 9614
rect 35196 9044 35252 9054
rect 35084 9042 35252 9044
rect 35084 8990 35198 9042
rect 35250 8990 35252 9042
rect 35084 8988 35252 8990
rect 35196 8978 35252 8988
rect 35420 9044 35476 9054
rect 35532 9044 35588 9548
rect 35644 9268 35700 10332
rect 35644 9174 35700 9212
rect 35420 9042 35588 9044
rect 35420 8990 35422 9042
rect 35474 8990 35588 9042
rect 35420 8988 35588 8990
rect 35420 8978 35476 8988
rect 35308 8930 35364 8942
rect 35308 8878 35310 8930
rect 35362 8878 35364 8930
rect 35308 8820 35364 8878
rect 34748 8764 35364 8820
rect 34748 8146 34804 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35420 8372 35476 8382
rect 34748 8094 34750 8146
rect 34802 8094 34804 8146
rect 34748 8082 34804 8094
rect 34972 8148 35028 8158
rect 34972 8054 35028 8092
rect 35420 8146 35476 8316
rect 35532 8260 35588 8988
rect 35756 8372 35812 10668
rect 35868 10610 35924 10780
rect 35980 10724 36036 12126
rect 36428 11620 36484 12460
rect 36428 11554 36484 11564
rect 36204 10724 36260 10734
rect 35980 10668 36204 10724
rect 35868 10558 35870 10610
rect 35922 10558 35924 10610
rect 35868 10546 35924 10558
rect 36204 10610 36260 10668
rect 36204 10558 36206 10610
rect 36258 10558 36260 10610
rect 36204 10546 36260 10558
rect 36428 10722 36484 10734
rect 36428 10670 36430 10722
rect 36482 10670 36484 10722
rect 35980 10500 36036 10510
rect 35980 10406 36036 10444
rect 36204 10164 36260 10174
rect 36204 9828 36260 10108
rect 36204 9826 36372 9828
rect 36204 9774 36206 9826
rect 36258 9774 36372 9826
rect 36204 9772 36372 9774
rect 36204 9762 36260 9772
rect 36092 9714 36148 9726
rect 36092 9662 36094 9714
rect 36146 9662 36148 9714
rect 35868 9602 35924 9614
rect 35868 9550 35870 9602
rect 35922 9550 35924 9602
rect 35868 9156 35924 9550
rect 35980 9604 36036 9614
rect 36092 9604 36148 9662
rect 36036 9548 36148 9604
rect 35980 9538 36036 9548
rect 35868 9062 35924 9100
rect 36316 9044 36372 9772
rect 36428 9268 36484 10670
rect 36764 10724 36820 10734
rect 36764 10630 36820 10668
rect 36428 9174 36484 9212
rect 36876 9268 36932 9278
rect 36876 9154 36932 9212
rect 36876 9102 36878 9154
rect 36930 9102 36932 9154
rect 36876 9090 36932 9102
rect 36652 9044 36708 9054
rect 35756 8306 35812 8316
rect 35980 9042 36372 9044
rect 35980 8990 36318 9042
rect 36370 8990 36372 9042
rect 35980 8988 36372 8990
rect 35644 8260 35700 8270
rect 35532 8204 35644 8260
rect 35644 8166 35700 8204
rect 35868 8260 35924 8270
rect 35980 8260 36036 8988
rect 36316 8978 36372 8988
rect 36540 9042 36708 9044
rect 36540 8990 36654 9042
rect 36706 8990 36708 9042
rect 36540 8988 36708 8990
rect 36316 8372 36372 8382
rect 36316 8278 36372 8316
rect 35868 8258 36036 8260
rect 35868 8206 35870 8258
rect 35922 8206 36036 8258
rect 35868 8204 36036 8206
rect 35868 8194 35924 8204
rect 35420 8094 35422 8146
rect 35474 8094 35476 8146
rect 35420 8082 35476 8094
rect 35756 8148 35812 8158
rect 35756 8054 35812 8092
rect 36540 8148 36596 8988
rect 36652 8978 36708 8988
rect 36764 8820 36820 8830
rect 36540 8082 36596 8092
rect 36652 8818 36820 8820
rect 36652 8766 36766 8818
rect 36818 8766 36820 8818
rect 36652 8764 36820 8766
rect 34188 7634 34244 7644
rect 34860 8034 34916 8046
rect 34860 7982 34862 8034
rect 34914 7982 34916 8034
rect 33516 6638 33518 6690
rect 33570 6638 33572 6690
rect 33516 6626 33572 6638
rect 31388 6526 31390 6578
rect 31442 6526 31444 6578
rect 31388 6514 31444 6526
rect 33404 6578 33460 6590
rect 33404 6526 33406 6578
rect 33458 6526 33460 6578
rect 32508 6468 32564 6478
rect 31276 5058 31332 5068
rect 32284 6466 32564 6468
rect 32284 6414 32510 6466
rect 32562 6414 32564 6466
rect 32284 6412 32564 6414
rect 31948 5010 32004 5022
rect 31948 4958 31950 5010
rect 32002 4958 32004 5010
rect 31948 4562 32004 4958
rect 31948 4510 31950 4562
rect 32002 4510 32004 4562
rect 31948 4498 32004 4510
rect 32284 4450 32340 6412
rect 32508 6402 32564 6412
rect 33404 5236 33460 6526
rect 34188 6466 34244 6478
rect 34188 6414 34190 6466
rect 34242 6414 34244 6466
rect 33404 5170 33460 5180
rect 33964 5906 34020 5918
rect 33964 5854 33966 5906
rect 34018 5854 34020 5906
rect 33964 5012 34020 5854
rect 34076 5236 34132 5246
rect 34188 5236 34244 6414
rect 34748 6020 34804 6030
rect 34860 6020 34916 7982
rect 36092 7588 36148 7598
rect 36316 7588 36372 7598
rect 36148 7586 36372 7588
rect 36148 7534 36318 7586
rect 36370 7534 36372 7586
rect 36148 7532 36372 7534
rect 36092 7494 36148 7532
rect 36316 7522 36372 7532
rect 36652 7474 36708 8764
rect 36764 8754 36820 8764
rect 37212 8260 37268 19294
rect 37884 19292 38276 19348
rect 37548 19236 37604 19246
rect 37884 19236 37940 19292
rect 38780 19236 38836 23436
rect 39228 23044 39284 27020
rect 39340 27412 39396 27422
rect 39340 26962 39396 27356
rect 39340 26910 39342 26962
rect 39394 26910 39396 26962
rect 39340 26898 39396 26910
rect 39340 24612 39396 24622
rect 39564 24612 39620 28028
rect 40012 28084 40068 29036
rect 40236 28644 40292 29484
rect 40348 29538 40404 29932
rect 40572 29894 40628 29932
rect 40348 29486 40350 29538
rect 40402 29486 40404 29538
rect 40348 29474 40404 29486
rect 40460 29428 40516 29438
rect 40236 28588 40404 28644
rect 40012 28018 40068 28028
rect 40124 28530 40180 28542
rect 40124 28478 40126 28530
rect 40178 28478 40180 28530
rect 40124 27860 40180 28478
rect 40236 28420 40292 28430
rect 40236 28326 40292 28364
rect 40236 28084 40292 28094
rect 40348 28084 40404 28588
rect 40460 28642 40516 29372
rect 40796 29426 40852 29438
rect 40796 29374 40798 29426
rect 40850 29374 40852 29426
rect 40796 28866 40852 29374
rect 40908 29204 40964 31388
rect 41132 29650 41188 31612
rect 41132 29598 41134 29650
rect 41186 29598 41188 29650
rect 41132 29586 41188 29598
rect 41132 29428 41188 29438
rect 41132 29334 41188 29372
rect 40908 29148 41188 29204
rect 40796 28814 40798 28866
rect 40850 28814 40852 28866
rect 40796 28802 40852 28814
rect 40460 28590 40462 28642
rect 40514 28590 40516 28642
rect 40460 28578 40516 28590
rect 40572 28644 40628 28654
rect 40460 28084 40516 28094
rect 40348 28082 40516 28084
rect 40348 28030 40462 28082
rect 40514 28030 40516 28082
rect 40348 28028 40516 28030
rect 40236 27990 40292 28028
rect 40460 28018 40516 28028
rect 39900 27858 40180 27860
rect 39900 27806 40126 27858
rect 40178 27806 40180 27858
rect 39900 27804 40180 27806
rect 39676 27412 39732 27422
rect 39676 26290 39732 27356
rect 39900 26516 39956 27804
rect 40124 27794 40180 27804
rect 40236 27524 40292 27534
rect 40236 27076 40292 27468
rect 40236 27074 40404 27076
rect 40236 27022 40238 27074
rect 40290 27022 40404 27074
rect 40236 27020 40404 27022
rect 40236 27010 40292 27020
rect 40012 26964 40068 27002
rect 40012 26898 40068 26908
rect 40348 26964 40404 27020
rect 40348 26898 40404 26908
rect 40124 26852 40180 26862
rect 40124 26850 40292 26852
rect 40124 26798 40126 26850
rect 40178 26798 40292 26850
rect 40124 26796 40292 26798
rect 40124 26786 40180 26796
rect 39900 26450 39956 26460
rect 40012 26628 40068 26638
rect 39676 26238 39678 26290
rect 39730 26238 39732 26290
rect 39676 25172 39732 26238
rect 39900 26180 39956 26190
rect 39900 26086 39956 26124
rect 40012 25956 40068 26572
rect 39676 25106 39732 25116
rect 39900 25900 40068 25956
rect 40124 26290 40180 26302
rect 40124 26238 40126 26290
rect 40178 26238 40180 26290
rect 39788 24612 39844 24622
rect 39564 24610 39844 24612
rect 39564 24558 39790 24610
rect 39842 24558 39844 24610
rect 39564 24556 39844 24558
rect 39340 24518 39396 24556
rect 39788 23492 39844 24556
rect 39788 23426 39844 23436
rect 39452 23268 39508 23278
rect 39452 23174 39508 23212
rect 39340 23044 39396 23054
rect 39228 23042 39396 23044
rect 39228 22990 39342 23042
rect 39394 22990 39396 23042
rect 39228 22988 39396 22990
rect 39340 22978 39396 22988
rect 39116 22932 39172 22942
rect 39116 22370 39172 22876
rect 39676 22932 39732 22942
rect 39676 22838 39732 22876
rect 39116 22318 39118 22370
rect 39170 22318 39172 22370
rect 39116 22306 39172 22318
rect 39788 21812 39844 21822
rect 39788 21698 39844 21756
rect 39788 21646 39790 21698
rect 39842 21646 39844 21698
rect 39788 21634 39844 21646
rect 39116 20804 39172 20814
rect 39116 20710 39172 20748
rect 39900 20244 39956 25900
rect 39900 20178 39956 20188
rect 40012 23604 40068 23614
rect 37548 19234 37940 19236
rect 37548 19182 37550 19234
rect 37602 19182 37940 19234
rect 37548 19180 37940 19182
rect 38668 19180 38836 19236
rect 39228 20132 39284 20142
rect 39228 19346 39284 20076
rect 39228 19294 39230 19346
rect 39282 19294 39284 19346
rect 37548 19170 37604 19180
rect 37996 19122 38052 19134
rect 37996 19070 37998 19122
rect 38050 19070 38052 19122
rect 37996 18564 38052 19070
rect 38108 18564 38164 18574
rect 37996 18562 38164 18564
rect 37996 18510 38110 18562
rect 38162 18510 38164 18562
rect 37996 18508 38164 18510
rect 38108 18498 38164 18508
rect 38444 18452 38500 18462
rect 38220 18450 38500 18452
rect 38220 18398 38446 18450
rect 38498 18398 38500 18450
rect 38220 18396 38500 18398
rect 37436 18338 37492 18350
rect 37436 18286 37438 18338
rect 37490 18286 37492 18338
rect 37324 15316 37380 15326
rect 37324 15222 37380 15260
rect 37436 12964 37492 18286
rect 37772 18340 37828 18350
rect 38220 18340 38276 18396
rect 38444 18386 38500 18396
rect 37772 18338 38276 18340
rect 37772 18286 37774 18338
rect 37826 18286 38276 18338
rect 37772 18284 38276 18286
rect 37772 18274 37828 18284
rect 38444 18226 38500 18238
rect 38444 18174 38446 18226
rect 38498 18174 38500 18226
rect 38220 17556 38276 17566
rect 37548 17444 37604 17454
rect 37548 16098 37604 17388
rect 38108 17442 38164 17454
rect 38108 17390 38110 17442
rect 38162 17390 38164 17442
rect 37996 17108 38052 17118
rect 37996 17014 38052 17052
rect 38108 16884 38164 17390
rect 38108 16818 38164 16828
rect 37548 16046 37550 16098
rect 37602 16046 37604 16098
rect 37548 16034 37604 16046
rect 37660 15876 37716 15886
rect 37660 15782 37716 15820
rect 38220 14532 38276 17500
rect 37548 13188 37604 13198
rect 37884 13188 37940 13198
rect 37604 13186 37940 13188
rect 37604 13134 37886 13186
rect 37938 13134 37940 13186
rect 37604 13132 37940 13134
rect 37548 13074 37604 13132
rect 37548 13022 37550 13074
rect 37602 13022 37604 13074
rect 37548 13010 37604 13022
rect 37436 12898 37492 12908
rect 37772 11954 37828 11966
rect 37772 11902 37774 11954
rect 37826 11902 37828 11954
rect 37324 11732 37380 11742
rect 37324 10836 37380 11676
rect 37324 10742 37380 10780
rect 37772 10164 37828 11902
rect 37884 11956 37940 13132
rect 38220 12962 38276 14476
rect 38332 16548 38388 16558
rect 38332 13748 38388 16492
rect 38444 16324 38500 18174
rect 38556 17444 38612 17454
rect 38556 17108 38612 17388
rect 38668 17220 38724 19180
rect 38780 19012 38836 19022
rect 39228 19012 39284 19294
rect 38836 18956 39284 19012
rect 39452 20020 39508 20030
rect 38780 18918 38836 18956
rect 39116 18562 39172 18574
rect 39116 18510 39118 18562
rect 39170 18510 39172 18562
rect 38892 18450 38948 18462
rect 38892 18398 38894 18450
rect 38946 18398 38948 18450
rect 38892 17892 38948 18398
rect 38892 17826 38948 17836
rect 38668 17154 38724 17164
rect 39004 17668 39060 17678
rect 38556 17042 38612 17052
rect 38668 16996 38724 17006
rect 38556 16884 38612 16894
rect 38668 16884 38724 16940
rect 38556 16882 38724 16884
rect 38556 16830 38558 16882
rect 38610 16830 38724 16882
rect 38556 16828 38724 16830
rect 38780 16882 38836 16894
rect 38780 16830 38782 16882
rect 38834 16830 38836 16882
rect 38556 16818 38612 16828
rect 38444 16268 38724 16324
rect 38556 15986 38612 15998
rect 38556 15934 38558 15986
rect 38610 15934 38612 15986
rect 38444 15874 38500 15886
rect 38444 15822 38446 15874
rect 38498 15822 38500 15874
rect 38444 14420 38500 15822
rect 38556 15764 38612 15934
rect 38556 15698 38612 15708
rect 38668 15148 38724 16268
rect 38780 15988 38836 16830
rect 39004 16884 39060 17612
rect 39004 16818 39060 16828
rect 39004 16100 39060 16110
rect 39004 16006 39060 16044
rect 38780 15932 38948 15988
rect 38780 15428 38836 15438
rect 38780 15334 38836 15372
rect 38668 15092 38836 15148
rect 38444 14354 38500 14364
rect 38780 14418 38836 15092
rect 38780 14366 38782 14418
rect 38834 14366 38836 14418
rect 38780 14354 38836 14366
rect 38556 13748 38612 13758
rect 38332 13746 38612 13748
rect 38332 13694 38558 13746
rect 38610 13694 38612 13746
rect 38332 13692 38612 13694
rect 38220 12910 38222 12962
rect 38274 12910 38276 12962
rect 38220 12898 38276 12910
rect 38332 12964 38388 12974
rect 37996 12738 38052 12750
rect 37996 12686 37998 12738
rect 38050 12686 38052 12738
rect 37996 12292 38052 12686
rect 37996 12226 38052 12236
rect 38108 12740 38164 12750
rect 38108 12180 38164 12684
rect 38108 12086 38164 12124
rect 38332 12178 38388 12908
rect 38332 12126 38334 12178
rect 38386 12126 38388 12178
rect 38332 12114 38388 12126
rect 37884 11890 37940 11900
rect 38556 10164 38612 13692
rect 38668 13522 38724 13534
rect 38668 13470 38670 13522
rect 38722 13470 38724 13522
rect 38668 13188 38724 13470
rect 38892 13188 38948 15932
rect 39116 15148 39172 18510
rect 39228 17556 39284 17566
rect 39228 17462 39284 17500
rect 39228 16996 39284 17006
rect 39452 16996 39508 19964
rect 39788 20020 39844 20030
rect 40012 20020 40068 23548
rect 39844 20018 40068 20020
rect 39844 19966 40014 20018
rect 40066 19966 40068 20018
rect 39844 19964 40068 19966
rect 39788 19926 39844 19964
rect 40012 19954 40068 19964
rect 40124 20130 40180 26238
rect 40236 26290 40292 26796
rect 40236 26238 40238 26290
rect 40290 26238 40292 26290
rect 40236 26226 40292 26238
rect 40348 24724 40404 24734
rect 40348 24630 40404 24668
rect 40572 23940 40628 28588
rect 40684 28530 40740 28542
rect 40684 28478 40686 28530
rect 40738 28478 40740 28530
rect 40684 27412 40740 28478
rect 40684 27346 40740 27356
rect 40796 28532 40852 28542
rect 40796 28418 40852 28476
rect 40796 28366 40798 28418
rect 40850 28366 40852 28418
rect 40684 27076 40740 27114
rect 40684 27010 40740 27020
rect 40796 26908 40852 28366
rect 41020 28420 41076 28430
rect 41020 28084 41076 28364
rect 41020 27990 41076 28028
rect 41132 27860 41188 29148
rect 40348 23884 40628 23940
rect 40684 26852 40852 26908
rect 40908 27804 41188 27860
rect 40236 21586 40292 21598
rect 40236 21534 40238 21586
rect 40290 21534 40292 21586
rect 40236 20804 40292 21534
rect 40236 20738 40292 20748
rect 40124 20078 40126 20130
rect 40178 20078 40180 20130
rect 39564 19124 39620 19134
rect 39564 19030 39620 19068
rect 40124 18562 40180 20078
rect 40124 18510 40126 18562
rect 40178 18510 40180 18562
rect 40124 18498 40180 18510
rect 39788 18452 39844 18462
rect 39676 18450 39844 18452
rect 39676 18398 39790 18450
rect 39842 18398 39844 18450
rect 39676 18396 39844 18398
rect 39564 17666 39620 17678
rect 39564 17614 39566 17666
rect 39618 17614 39620 17666
rect 39564 17444 39620 17614
rect 39564 17378 39620 17388
rect 39676 17108 39732 18396
rect 39788 18386 39844 18396
rect 40348 18452 40404 23884
rect 40572 22258 40628 22270
rect 40572 22206 40574 22258
rect 40626 22206 40628 22258
rect 40572 21588 40628 22206
rect 40572 20690 40628 21532
rect 40572 20638 40574 20690
rect 40626 20638 40628 20690
rect 40572 20626 40628 20638
rect 40684 19236 40740 26852
rect 40908 26178 40964 27804
rect 41020 26964 41076 27002
rect 41020 26898 41076 26908
rect 40908 26126 40910 26178
rect 40962 26126 40964 26178
rect 40796 25284 40852 25294
rect 40796 24050 40852 25228
rect 40796 23998 40798 24050
rect 40850 23998 40852 24050
rect 40796 23986 40852 23998
rect 40908 23604 40964 26126
rect 41244 24948 41300 32732
rect 42252 32722 42308 32734
rect 41804 32564 41860 32574
rect 41804 32470 41860 32508
rect 42028 32562 42084 32574
rect 42364 32564 42420 34412
rect 42700 34690 42868 34692
rect 42700 34638 42814 34690
rect 42866 34638 42868 34690
rect 42700 34636 42868 34638
rect 42588 34020 42644 34030
rect 42588 33926 42644 33964
rect 42588 33684 42644 33694
rect 42476 33124 42532 33134
rect 42476 32674 42532 33068
rect 42588 32786 42644 33628
rect 42700 33346 42756 34636
rect 42812 34626 42868 34636
rect 43372 34690 43428 35196
rect 43372 34638 43374 34690
rect 43426 34638 43428 34690
rect 42924 34242 42980 34254
rect 42924 34190 42926 34242
rect 42978 34190 42980 34242
rect 42924 34020 42980 34190
rect 42924 33954 42980 33964
rect 43036 34130 43092 34142
rect 43036 34078 43038 34130
rect 43090 34078 43092 34130
rect 42700 33294 42702 33346
rect 42754 33294 42756 33346
rect 42700 33282 42756 33294
rect 43036 33124 43092 34078
rect 43036 33058 43092 33068
rect 43148 33346 43204 33358
rect 43148 33294 43150 33346
rect 43202 33294 43204 33346
rect 43148 32900 43204 33294
rect 43372 33348 43428 34638
rect 43708 35140 43764 35150
rect 44044 35140 44100 36206
rect 44156 36204 44268 36260
rect 44156 35922 44212 36204
rect 44268 36194 44324 36204
rect 44156 35870 44158 35922
rect 44210 35870 44212 35922
rect 44156 35858 44212 35870
rect 44380 35922 44436 37660
rect 44380 35870 44382 35922
rect 44434 35870 44436 35922
rect 44380 35858 44436 35870
rect 44268 35812 44324 35822
rect 44268 35700 44324 35756
rect 44380 35700 44436 35710
rect 44268 35698 44436 35700
rect 44268 35646 44382 35698
rect 44434 35646 44436 35698
rect 44268 35644 44436 35646
rect 44380 35634 44436 35644
rect 43484 33572 43540 33582
rect 43484 33478 43540 33516
rect 43372 33292 43540 33348
rect 43148 32834 43204 32844
rect 42588 32734 42590 32786
rect 42642 32734 42644 32786
rect 42588 32722 42644 32734
rect 42476 32622 42478 32674
rect 42530 32622 42532 32674
rect 42476 32610 42532 32622
rect 42028 32510 42030 32562
rect 42082 32510 42084 32562
rect 42028 32116 42084 32510
rect 42028 32050 42084 32060
rect 42252 32508 42420 32564
rect 43260 32564 43316 32574
rect 42140 31108 42196 31118
rect 42140 30324 42196 31052
rect 42140 30210 42196 30268
rect 42140 30158 42142 30210
rect 42194 30158 42196 30210
rect 42140 30146 42196 30158
rect 41356 29988 41412 29998
rect 41356 29426 41412 29932
rect 41356 29374 41358 29426
rect 41410 29374 41412 29426
rect 41356 29362 41412 29374
rect 42028 29652 42084 29662
rect 42028 29426 42084 29596
rect 42028 29374 42030 29426
rect 42082 29374 42084 29426
rect 42028 29362 42084 29374
rect 41356 28644 41412 28654
rect 41356 28550 41412 28588
rect 41804 28532 41860 28542
rect 41804 28438 41860 28476
rect 41468 27748 41524 27758
rect 41468 27076 41524 27692
rect 41468 26982 41524 27020
rect 42252 26908 42308 32508
rect 43260 32450 43316 32508
rect 43260 32398 43262 32450
rect 43314 32398 43316 32450
rect 42812 31556 42868 31566
rect 42588 30212 42644 30222
rect 42588 29986 42644 30156
rect 42588 29934 42590 29986
rect 42642 29934 42644 29986
rect 42588 28868 42644 29934
rect 42700 29316 42756 29326
rect 42700 29222 42756 29260
rect 42588 28802 42644 28812
rect 42700 28532 42756 28542
rect 42812 28532 42868 31500
rect 43148 30212 43204 30222
rect 43148 30118 43204 30156
rect 42756 28476 42868 28532
rect 43148 29988 43204 29998
rect 42700 28466 42756 28476
rect 42252 26852 42532 26908
rect 41244 24882 41300 24892
rect 42476 24946 42532 26852
rect 43036 26180 43092 26190
rect 43036 26086 43092 26124
rect 42476 24894 42478 24946
rect 42530 24894 42532 24946
rect 42476 24882 42532 24894
rect 40908 23538 40964 23548
rect 41244 24724 41300 24734
rect 41244 23378 41300 24668
rect 42700 24722 42756 24734
rect 42700 24670 42702 24722
rect 42754 24670 42756 24722
rect 42364 24610 42420 24622
rect 42364 24558 42366 24610
rect 42418 24558 42420 24610
rect 41244 23326 41246 23378
rect 41298 23326 41300 23378
rect 41244 23314 41300 23326
rect 41356 23938 41412 23950
rect 41356 23886 41358 23938
rect 41410 23886 41412 23938
rect 41356 23268 41412 23886
rect 42140 23828 42196 23838
rect 42364 23828 42420 24558
rect 42140 23826 42420 23828
rect 42140 23774 42142 23826
rect 42194 23774 42420 23826
rect 42140 23772 42420 23774
rect 41804 23268 41860 23278
rect 41244 23154 41300 23166
rect 41244 23102 41246 23154
rect 41298 23102 41300 23154
rect 41244 22820 41300 23102
rect 41244 22754 41300 22764
rect 41132 22370 41188 22382
rect 41132 22318 41134 22370
rect 41186 22318 41188 22370
rect 41020 21364 41076 21374
rect 41020 21270 41076 21308
rect 41020 21140 41076 21150
rect 41020 19908 41076 21084
rect 41132 20132 41188 22318
rect 41356 21588 41412 23212
rect 41580 23212 41804 23268
rect 41580 23154 41636 23212
rect 41804 23202 41860 23212
rect 41580 23102 41582 23154
rect 41634 23102 41636 23154
rect 41580 23090 41636 23102
rect 42028 23156 42084 23166
rect 42140 23156 42196 23772
rect 42700 23268 42756 24670
rect 42700 23202 42756 23212
rect 42924 24722 42980 24734
rect 42924 24670 42926 24722
rect 42978 24670 42980 24722
rect 42924 23940 42980 24670
rect 43036 23940 43092 23950
rect 42924 23938 43092 23940
rect 42924 23886 43038 23938
rect 43090 23886 43092 23938
rect 42924 23884 43092 23886
rect 42028 23154 42196 23156
rect 42028 23102 42030 23154
rect 42082 23102 42196 23154
rect 42028 23100 42196 23102
rect 42028 23090 42084 23100
rect 42140 23044 42196 23100
rect 42140 22978 42196 22988
rect 42588 23042 42644 23054
rect 42588 22990 42590 23042
rect 42642 22990 42644 23042
rect 41804 22932 41860 22942
rect 41804 22482 41860 22876
rect 41804 22430 41806 22482
rect 41858 22430 41860 22482
rect 41580 22148 41636 22158
rect 41580 22054 41636 22092
rect 41580 21588 41636 21598
rect 41356 21532 41580 21588
rect 41580 21494 41636 21532
rect 41804 21586 41860 22430
rect 42588 22932 42644 22990
rect 42476 22370 42532 22382
rect 42476 22318 42478 22370
rect 42530 22318 42532 22370
rect 42140 22258 42196 22270
rect 42140 22206 42142 22258
rect 42194 22206 42196 22258
rect 42140 21812 42196 22206
rect 42476 22036 42532 22318
rect 42476 21970 42532 21980
rect 42140 21746 42196 21756
rect 42364 21700 42420 21710
rect 42364 21606 42420 21644
rect 41804 21534 41806 21586
rect 41858 21534 41860 21586
rect 41244 21476 41300 21486
rect 41244 21474 41412 21476
rect 41244 21422 41246 21474
rect 41298 21422 41412 21474
rect 41244 21420 41412 21422
rect 41244 21410 41300 21420
rect 41132 20066 41188 20076
rect 41020 19906 41188 19908
rect 41020 19854 41022 19906
rect 41074 19854 41188 19906
rect 41020 19852 41188 19854
rect 41020 19842 41076 19852
rect 40348 18386 40404 18396
rect 40460 19180 40740 19236
rect 40236 18338 40292 18350
rect 40236 18286 40238 18338
rect 40290 18286 40292 18338
rect 40236 17220 40292 18286
rect 40236 17154 40292 17164
rect 39228 16994 39508 16996
rect 39228 16942 39230 16994
rect 39282 16942 39508 16994
rect 39228 16940 39508 16942
rect 39228 16930 39284 16940
rect 39452 16884 39508 16940
rect 39452 16818 39508 16828
rect 39564 17052 39732 17108
rect 39228 16770 39284 16782
rect 39228 16718 39230 16770
rect 39282 16718 39284 16770
rect 39228 15988 39284 16718
rect 39228 15922 39284 15932
rect 39340 16772 39396 16782
rect 39004 15092 39172 15148
rect 39228 15538 39284 15550
rect 39228 15486 39230 15538
rect 39282 15486 39284 15538
rect 39004 13860 39060 15092
rect 39228 14530 39284 15486
rect 39340 15314 39396 16716
rect 39564 16548 39620 17052
rect 40012 16996 40068 17006
rect 39564 16482 39620 16492
rect 39676 16994 40068 16996
rect 39676 16942 40014 16994
rect 40066 16942 40068 16994
rect 39676 16940 40068 16942
rect 39676 16212 39732 16940
rect 40012 16930 40068 16940
rect 40236 16996 40292 17006
rect 40460 16996 40516 19180
rect 40572 19010 40628 19022
rect 40572 18958 40574 19010
rect 40626 18958 40628 19010
rect 40572 17668 40628 18958
rect 41132 18564 41188 19852
rect 41244 19236 41300 19246
rect 41244 19142 41300 19180
rect 41356 19124 41412 21420
rect 41468 20916 41524 20926
rect 41468 20802 41524 20860
rect 41468 20750 41470 20802
rect 41522 20750 41524 20802
rect 41468 20738 41524 20750
rect 41580 20692 41636 20702
rect 41580 20578 41636 20636
rect 41580 20526 41582 20578
rect 41634 20526 41636 20578
rect 41580 20514 41636 20526
rect 41692 20580 41748 20590
rect 41692 20486 41748 20524
rect 41804 20356 41860 21534
rect 41692 20300 41860 20356
rect 42028 21028 42084 21038
rect 42028 20914 42084 20972
rect 42028 20862 42030 20914
rect 42082 20862 42084 20914
rect 41580 20132 41636 20142
rect 41468 20020 41524 20030
rect 41468 19926 41524 19964
rect 41356 19058 41412 19068
rect 41580 19234 41636 20076
rect 41580 19182 41582 19234
rect 41634 19182 41636 19234
rect 41244 18564 41300 18574
rect 41132 18562 41300 18564
rect 41132 18510 41246 18562
rect 41298 18510 41300 18562
rect 41132 18508 41300 18510
rect 41244 18498 41300 18508
rect 40908 18452 40964 18462
rect 40684 17780 40740 17790
rect 40684 17686 40740 17724
rect 40572 17602 40628 17612
rect 40292 16940 40516 16996
rect 39340 15262 39342 15314
rect 39394 15262 39396 15314
rect 39340 15250 39396 15262
rect 39452 16156 39732 16212
rect 40236 16882 40292 16940
rect 40236 16830 40238 16882
rect 40290 16830 40292 16882
rect 40236 16212 40292 16830
rect 39452 16098 39508 16156
rect 39452 16046 39454 16098
rect 39506 16046 39508 16098
rect 39452 15148 39508 16046
rect 40236 16098 40292 16156
rect 40236 16046 40238 16098
rect 40290 16046 40292 16098
rect 40236 16034 40292 16046
rect 40348 16324 40404 16334
rect 39788 15988 39844 15998
rect 39228 14478 39230 14530
rect 39282 14478 39284 14530
rect 39228 14466 39284 14478
rect 39340 15092 39508 15148
rect 39564 15876 39620 15886
rect 39004 13794 39060 13804
rect 39340 13858 39396 15092
rect 39340 13806 39342 13858
rect 39394 13806 39396 13858
rect 39340 13794 39396 13806
rect 38668 13132 38948 13188
rect 38668 12964 38724 12974
rect 38668 12962 38836 12964
rect 38668 12910 38670 12962
rect 38722 12910 38836 12962
rect 38668 12908 38836 12910
rect 38668 12898 38724 12908
rect 38668 12404 38724 12414
rect 38668 12310 38724 12348
rect 38780 12180 38836 12908
rect 38780 12114 38836 12124
rect 38780 10724 38836 10734
rect 38780 10610 38836 10668
rect 38780 10558 38782 10610
rect 38834 10558 38836 10610
rect 38780 10546 38836 10558
rect 37772 10098 37828 10108
rect 38220 10108 38612 10164
rect 38108 9156 38164 9166
rect 38108 9062 38164 9100
rect 37100 8258 37268 8260
rect 37100 8206 37214 8258
rect 37266 8206 37268 8258
rect 37100 8204 37268 8206
rect 36988 8148 37044 8158
rect 36988 8054 37044 8092
rect 36652 7422 36654 7474
rect 36706 7422 36708 7474
rect 36652 7410 36708 7422
rect 36988 7476 37044 7486
rect 36988 7382 37044 7420
rect 36764 7362 36820 7374
rect 36764 7310 36766 7362
rect 36818 7310 36820 7362
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34748 6018 34916 6020
rect 34748 5966 34750 6018
rect 34802 5966 34916 6018
rect 34748 5964 34916 5966
rect 34748 5954 34804 5964
rect 36764 5796 36820 7310
rect 37100 6692 37156 8204
rect 37212 8194 37268 8204
rect 37884 7588 37940 7598
rect 37884 7494 37940 7532
rect 38220 7586 38276 10108
rect 38892 10052 38948 13132
rect 39116 13746 39172 13758
rect 39116 13694 39118 13746
rect 39170 13694 39172 13746
rect 39116 13636 39172 13694
rect 39116 12964 39172 13580
rect 39564 13076 39620 15820
rect 39788 14530 39844 15932
rect 40348 15764 40404 16268
rect 40236 15540 40292 15550
rect 40348 15540 40404 15708
rect 40236 15538 40404 15540
rect 40236 15486 40238 15538
rect 40290 15486 40404 15538
rect 40236 15484 40404 15486
rect 40236 15474 40292 15484
rect 39788 14478 39790 14530
rect 39842 14478 39844 14530
rect 39788 14466 39844 14478
rect 40796 14642 40852 14654
rect 40796 14590 40798 14642
rect 40850 14590 40852 14642
rect 39676 14420 39732 14430
rect 40124 14420 40180 14430
rect 39676 14326 39732 14364
rect 40012 14364 40124 14420
rect 40012 13970 40068 14364
rect 40124 14354 40180 14364
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 40012 13906 40068 13918
rect 40124 13860 40180 13870
rect 40124 13766 40180 13804
rect 39676 13748 39732 13758
rect 39676 13654 39732 13692
rect 39900 13746 39956 13758
rect 39900 13694 39902 13746
rect 39954 13694 39956 13746
rect 39116 12870 39172 12908
rect 39340 13020 39620 13076
rect 39004 12290 39060 12302
rect 39004 12238 39006 12290
rect 39058 12238 39060 12290
rect 39004 12068 39060 12238
rect 39004 12002 39060 12012
rect 38332 9996 38948 10052
rect 39004 11844 39060 11854
rect 39004 10722 39060 11788
rect 39004 10670 39006 10722
rect 39058 10670 39060 10722
rect 38332 9268 38388 9996
rect 38332 9174 38388 9212
rect 38444 9826 38500 9838
rect 38444 9774 38446 9826
rect 38498 9774 38500 9826
rect 38444 8930 38500 9774
rect 38668 9828 38724 9838
rect 38668 9734 38724 9772
rect 38444 8878 38446 8930
rect 38498 8878 38500 8930
rect 38220 7534 38222 7586
rect 38274 7534 38276 7586
rect 37996 7476 38052 7486
rect 37996 7382 38052 7420
rect 36204 5740 36820 5796
rect 36876 6636 37156 6692
rect 36876 5794 36932 6636
rect 36876 5742 36878 5794
rect 36930 5742 36932 5794
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34132 5180 34244 5236
rect 34076 5142 34132 5180
rect 33964 4946 34020 4956
rect 35420 5012 35476 5022
rect 32284 4398 32286 4450
rect 32338 4398 32340 4450
rect 32284 4386 32340 4398
rect 30604 4338 31220 4340
rect 30604 4286 30606 4338
rect 30658 4286 31220 4338
rect 30604 4284 31220 4286
rect 35420 4338 35476 4956
rect 36204 4450 36260 5740
rect 36876 5730 36932 5742
rect 37324 5794 37380 5806
rect 37324 5742 37326 5794
rect 37378 5742 37380 5794
rect 37324 5012 37380 5742
rect 37324 4946 37380 4956
rect 37996 5122 38052 5134
rect 37996 5070 37998 5122
rect 38050 5070 38052 5122
rect 37996 5012 38052 5070
rect 37996 4946 38052 4956
rect 36204 4398 36206 4450
rect 36258 4398 36260 4450
rect 36204 4386 36260 4398
rect 35420 4286 35422 4338
rect 35474 4286 35476 4338
rect 27468 3668 27524 3678
rect 27244 3666 27524 3668
rect 27244 3614 27470 3666
rect 27522 3614 27524 3666
rect 27244 3612 27524 3614
rect 25340 3602 25396 3612
rect 27468 3602 27524 3612
rect 29820 3666 29876 3678
rect 29820 3614 29822 3666
rect 29874 3614 29876 3666
rect 29820 3388 29876 3614
rect 30604 3556 30660 4284
rect 35420 4274 35476 4286
rect 38220 4228 38276 7534
rect 38332 8596 38388 8606
rect 38332 7586 38388 8540
rect 38444 8428 38500 8878
rect 38892 9714 38948 9726
rect 38892 9662 38894 9714
rect 38946 9662 38948 9714
rect 38892 8596 38948 9662
rect 39004 9604 39060 10670
rect 39116 10500 39172 10510
rect 39116 9826 39172 10444
rect 39340 10164 39396 13020
rect 39564 12852 39620 12862
rect 39564 12758 39620 12796
rect 39900 11844 39956 13694
rect 40236 13746 40292 13758
rect 40236 13694 40238 13746
rect 40290 13694 40292 13746
rect 40236 13636 40292 13694
rect 40124 13580 40292 13636
rect 40124 12068 40180 13580
rect 40124 12002 40180 12012
rect 40236 13412 40292 13422
rect 39900 11778 39956 11788
rect 39452 10722 39508 10734
rect 39452 10670 39454 10722
rect 39506 10670 39508 10722
rect 39452 10500 39508 10670
rect 39564 10724 39620 10734
rect 39564 10630 39620 10668
rect 39452 10434 39508 10444
rect 39676 10386 39732 10398
rect 39676 10334 39678 10386
rect 39730 10334 39732 10386
rect 39676 10164 39732 10334
rect 39340 10108 39508 10164
rect 39228 10052 39284 10062
rect 39228 9958 39284 9996
rect 39116 9774 39118 9826
rect 39170 9774 39172 9826
rect 39116 9762 39172 9774
rect 39004 9548 39284 9604
rect 38892 8530 38948 8540
rect 38444 8372 38948 8428
rect 38892 8258 38948 8372
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38892 8194 38948 8206
rect 39228 8034 39284 9548
rect 39228 7982 39230 8034
rect 39282 7982 39284 8034
rect 39228 7924 39284 7982
rect 39228 7858 39284 7868
rect 39340 8370 39396 8382
rect 39340 8318 39342 8370
rect 39394 8318 39396 8370
rect 38780 7700 38836 7710
rect 38332 7534 38334 7586
rect 38386 7534 38388 7586
rect 38332 6692 38388 7534
rect 38668 7588 38724 7598
rect 38668 7494 38724 7532
rect 38332 6626 38388 6636
rect 38780 5234 38836 7644
rect 39004 7700 39060 7738
rect 39004 7634 39060 7644
rect 38892 7474 38948 7486
rect 38892 7422 38894 7474
rect 38946 7422 38948 7474
rect 38892 6916 38948 7422
rect 39340 7474 39396 8318
rect 39452 8146 39508 10108
rect 39676 10098 39732 10108
rect 39452 8094 39454 8146
rect 39506 8094 39508 8146
rect 39452 7588 39508 8094
rect 39564 7588 39620 7598
rect 39452 7586 39620 7588
rect 39452 7534 39566 7586
rect 39618 7534 39620 7586
rect 39452 7532 39620 7534
rect 39564 7522 39620 7532
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39340 7410 39396 7422
rect 39788 7474 39844 7486
rect 39788 7422 39790 7474
rect 39842 7422 39844 7474
rect 39228 6916 39284 6926
rect 38892 6914 39284 6916
rect 38892 6862 39230 6914
rect 39282 6862 39284 6914
rect 38892 6860 39284 6862
rect 39228 6850 39284 6860
rect 39116 6692 39172 6702
rect 39116 6598 39172 6636
rect 38780 5182 38782 5234
rect 38834 5182 38836 5234
rect 38780 5170 38836 5182
rect 39228 6468 39284 6478
rect 39788 6468 39844 7422
rect 39228 6466 39844 6468
rect 39228 6414 39230 6466
rect 39282 6414 39844 6466
rect 39228 6412 39844 6414
rect 39228 5236 39284 6412
rect 39228 5170 39284 5180
rect 38780 4340 38836 4350
rect 38780 4246 38836 4284
rect 38332 4228 38388 4238
rect 38220 4226 38388 4228
rect 38220 4174 38334 4226
rect 38386 4174 38388 4226
rect 38220 4172 38388 4174
rect 38332 4162 38388 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 30604 3490 30660 3500
rect 34076 3668 34132 3678
rect 29596 3332 29876 3388
rect 29596 800 29652 3332
rect 34076 800 34132 3612
rect 36988 3668 37044 3678
rect 36988 3574 37044 3612
rect 40236 3666 40292 13356
rect 40460 12852 40516 12862
rect 40460 12758 40516 12796
rect 40684 12738 40740 12750
rect 40684 12686 40686 12738
rect 40738 12686 40740 12738
rect 40684 11844 40740 12686
rect 40684 11778 40740 11788
rect 40796 11396 40852 14590
rect 40908 14644 40964 18396
rect 41468 18452 41524 18462
rect 41580 18452 41636 19182
rect 41468 18450 41636 18452
rect 41468 18398 41470 18450
rect 41522 18398 41636 18450
rect 41468 18396 41636 18398
rect 41692 19236 41748 20300
rect 41916 20244 41972 20254
rect 42028 20244 42084 20862
rect 41916 20242 42084 20244
rect 41916 20190 41918 20242
rect 41970 20190 42084 20242
rect 41916 20188 42084 20190
rect 42140 20804 42196 20814
rect 42140 20244 42196 20748
rect 42476 20802 42532 20814
rect 42476 20750 42478 20802
rect 42530 20750 42532 20802
rect 42252 20244 42308 20254
rect 42140 20242 42308 20244
rect 42140 20190 42254 20242
rect 42306 20190 42308 20242
rect 42140 20188 42308 20190
rect 41916 20178 41972 20188
rect 42252 20178 42308 20188
rect 42476 20244 42532 20750
rect 42476 20178 42532 20188
rect 41804 20132 41860 20142
rect 41804 20038 41860 20076
rect 41692 18450 41748 19180
rect 42140 20020 42196 20030
rect 41692 18398 41694 18450
rect 41746 18398 41748 18450
rect 41468 18386 41524 18396
rect 41692 18386 41748 18398
rect 41916 19124 41972 19134
rect 41916 18450 41972 19068
rect 42140 19124 42196 19964
rect 42364 19908 42420 19918
rect 42588 19908 42644 22876
rect 42700 21812 42756 21822
rect 42924 21812 42980 23884
rect 43036 23874 43092 23884
rect 43148 23380 43204 29932
rect 43260 26908 43316 32398
rect 43372 31780 43428 31790
rect 43372 31686 43428 31724
rect 43372 31444 43428 31454
rect 43484 31444 43540 33292
rect 43708 32786 43764 35084
rect 43820 35084 44100 35140
rect 44156 35588 44212 35598
rect 43820 34130 43876 35084
rect 44156 35028 44212 35532
rect 43820 34078 43822 34130
rect 43874 34078 43876 34130
rect 43820 34066 43876 34078
rect 44044 34972 44212 35028
rect 43708 32734 43710 32786
rect 43762 32734 43764 32786
rect 43708 32722 43764 32734
rect 43428 31388 43540 31444
rect 43596 32562 43652 32574
rect 43596 32510 43598 32562
rect 43650 32510 43652 32562
rect 43372 31378 43428 31388
rect 43372 30324 43428 30334
rect 43372 30210 43428 30268
rect 43596 30322 43652 32510
rect 43932 32562 43988 32574
rect 43932 32510 43934 32562
rect 43986 32510 43988 32562
rect 43932 32452 43988 32510
rect 43932 32386 43988 32396
rect 43820 31892 43876 31902
rect 43820 31220 43876 31836
rect 43820 31126 43876 31164
rect 43596 30270 43598 30322
rect 43650 30270 43652 30322
rect 43596 30258 43652 30270
rect 43372 30158 43374 30210
rect 43426 30158 43428 30210
rect 43372 30146 43428 30158
rect 43596 29988 43652 29998
rect 43484 29986 43652 29988
rect 43484 29934 43598 29986
rect 43650 29934 43652 29986
rect 43484 29932 43652 29934
rect 43484 28868 43540 29932
rect 43596 29922 43652 29932
rect 43708 29986 43764 29998
rect 43708 29934 43710 29986
rect 43762 29934 43764 29986
rect 43484 28802 43540 28812
rect 43708 27300 43764 29934
rect 43708 26908 43764 27244
rect 43260 26852 43428 26908
rect 43372 25284 43428 26852
rect 43372 25190 43428 25228
rect 43484 26852 43764 26908
rect 43820 29652 43876 29662
rect 43484 23380 43540 26852
rect 43820 26290 43876 29596
rect 43820 26238 43822 26290
rect 43874 26238 43876 26290
rect 43820 26180 43876 26238
rect 43820 26114 43876 26124
rect 43708 25508 43764 25518
rect 43708 24946 43764 25452
rect 44044 25396 44100 34972
rect 44380 34692 44436 34702
rect 44380 34598 44436 34636
rect 44380 34356 44436 34366
rect 44380 34242 44436 34300
rect 44380 34190 44382 34242
rect 44434 34190 44436 34242
rect 44380 34178 44436 34190
rect 44156 34132 44212 34142
rect 44156 34038 44212 34076
rect 44492 33572 44548 37884
rect 45164 37156 45220 38892
rect 45500 38724 45556 40350
rect 46060 39732 46116 43596
rect 46284 42084 46340 44046
rect 46732 43652 46788 43662
rect 46732 42868 46788 43596
rect 47292 43538 47348 45724
rect 47740 45714 47796 45724
rect 47852 45332 47908 46734
rect 48076 46676 48132 46686
rect 48076 46674 48244 46676
rect 48076 46622 48078 46674
rect 48130 46622 48244 46674
rect 48076 46620 48244 46622
rect 48076 46610 48132 46620
rect 47852 45266 47908 45276
rect 48076 46002 48132 46014
rect 48076 45950 48078 46002
rect 48130 45950 48132 46002
rect 48076 45330 48132 45950
rect 48188 45890 48244 46620
rect 48188 45838 48190 45890
rect 48242 45838 48244 45890
rect 48188 45826 48244 45838
rect 48300 46004 48356 48750
rect 48972 48356 49028 48972
rect 48972 48242 49028 48300
rect 48972 48190 48974 48242
rect 49026 48190 49028 48242
rect 48972 48178 49028 48190
rect 49084 49026 49252 49028
rect 49084 48974 49198 49026
rect 49250 48974 49252 49026
rect 49084 48972 49252 48974
rect 48748 48132 48804 48142
rect 48748 48130 48916 48132
rect 48748 48078 48750 48130
rect 48802 48078 48916 48130
rect 48748 48076 48916 48078
rect 48748 48066 48804 48076
rect 48860 48020 48916 48076
rect 49084 48020 49140 48972
rect 49196 48962 49252 48972
rect 49196 48132 49252 48142
rect 49196 48038 49252 48076
rect 48860 47964 49140 48020
rect 48748 47346 48804 47358
rect 48748 47294 48750 47346
rect 48802 47294 48804 47346
rect 48748 46340 48804 47294
rect 48860 47234 48916 47964
rect 49084 47572 49140 47582
rect 49084 47458 49140 47516
rect 49084 47406 49086 47458
rect 49138 47406 49140 47458
rect 49084 47394 49140 47406
rect 48860 47182 48862 47234
rect 48914 47182 48916 47234
rect 48860 46564 48916 47182
rect 49420 47124 49476 49756
rect 49980 49588 50036 49982
rect 51100 49924 51156 49934
rect 51324 49924 51380 51214
rect 51436 50596 51492 51326
rect 51660 51380 51716 51390
rect 51660 51286 51716 51324
rect 51436 50530 51492 50540
rect 51996 50594 52052 50606
rect 51996 50542 51998 50594
rect 52050 50542 52052 50594
rect 51100 49922 51380 49924
rect 51100 49870 51102 49922
rect 51154 49870 51380 49922
rect 51100 49868 51380 49870
rect 51100 49858 51156 49868
rect 49532 49532 50036 49588
rect 50428 49810 50484 49822
rect 50428 49758 50430 49810
rect 50482 49758 50484 49810
rect 49532 48468 49588 49532
rect 49644 49028 49700 49038
rect 49644 49026 49812 49028
rect 49644 48974 49646 49026
rect 49698 48974 49812 49026
rect 49644 48972 49812 48974
rect 49644 48962 49700 48972
rect 49644 48468 49700 48478
rect 49532 48466 49700 48468
rect 49532 48414 49646 48466
rect 49698 48414 49700 48466
rect 49532 48412 49700 48414
rect 49644 48402 49700 48412
rect 49644 47572 49700 47582
rect 49644 47478 49700 47516
rect 49532 47460 49588 47470
rect 49532 47366 49588 47404
rect 49420 47068 49588 47124
rect 48860 46498 48916 46508
rect 48748 46274 48804 46284
rect 48076 45278 48078 45330
rect 48130 45278 48132 45330
rect 48076 45266 48132 45278
rect 48188 45220 48244 45230
rect 48300 45220 48356 45948
rect 49196 46004 49252 46014
rect 49196 45890 49252 45948
rect 49196 45838 49198 45890
rect 49250 45838 49252 45890
rect 49196 45826 49252 45838
rect 49420 45890 49476 45902
rect 49420 45838 49422 45890
rect 49474 45838 49476 45890
rect 49084 45778 49140 45790
rect 49084 45726 49086 45778
rect 49138 45726 49140 45778
rect 49084 45556 49140 45726
rect 49084 45490 49140 45500
rect 48748 45332 48804 45342
rect 49420 45332 49476 45838
rect 48748 45238 48804 45276
rect 48860 45276 49476 45332
rect 48188 45218 48356 45220
rect 48188 45166 48190 45218
rect 48242 45166 48356 45218
rect 48188 45164 48356 45166
rect 48860 45218 48916 45276
rect 48860 45166 48862 45218
rect 48914 45166 48916 45218
rect 48188 45154 48244 45164
rect 47852 45106 47908 45118
rect 47852 45054 47854 45106
rect 47906 45054 47908 45106
rect 47516 44996 47572 45006
rect 47852 44996 47908 45054
rect 47516 44994 47908 44996
rect 47516 44942 47518 44994
rect 47570 44942 47908 44994
rect 47516 44940 47908 44942
rect 47516 44884 47572 44940
rect 47516 44818 47572 44828
rect 47516 44322 47572 44334
rect 47516 44270 47518 44322
rect 47570 44270 47572 44322
rect 47516 43764 47572 44270
rect 47740 44098 47796 44110
rect 47740 44046 47742 44098
rect 47794 44046 47796 44098
rect 47628 43764 47684 43774
rect 47516 43762 47684 43764
rect 47516 43710 47630 43762
rect 47682 43710 47684 43762
rect 47516 43708 47684 43710
rect 47628 43698 47684 43708
rect 47292 43486 47294 43538
rect 47346 43486 47348 43538
rect 47292 43474 47348 43486
rect 46844 43428 46900 43438
rect 47068 43428 47124 43438
rect 46844 43426 47236 43428
rect 46844 43374 46846 43426
rect 46898 43374 47070 43426
rect 47122 43374 47236 43426
rect 46844 43372 47236 43374
rect 46844 43362 46900 43372
rect 47068 43362 47124 43372
rect 46732 42866 47124 42868
rect 46732 42814 46734 42866
rect 46786 42814 47124 42866
rect 46732 42812 47124 42814
rect 46732 42802 46788 42812
rect 47068 42756 47124 42812
rect 47068 42662 47124 42700
rect 46284 42018 46340 42028
rect 46732 41860 46788 41870
rect 46732 41766 46788 41804
rect 47180 40628 47236 43372
rect 47740 42868 47796 44046
rect 48860 43316 48916 45166
rect 49532 43708 49588 47068
rect 49756 45780 49812 48972
rect 50428 47572 50484 49758
rect 51884 49138 51940 49150
rect 51884 49086 51886 49138
rect 51938 49086 51940 49138
rect 51884 48916 51940 49086
rect 51884 48850 51940 48860
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50316 47516 50484 47572
rect 50876 48242 50932 48254
rect 50876 48190 50878 48242
rect 50930 48190 50932 48242
rect 50316 47124 50372 47516
rect 50428 47348 50484 47358
rect 50764 47348 50820 47358
rect 50428 47346 50820 47348
rect 50428 47294 50430 47346
rect 50482 47294 50766 47346
rect 50818 47294 50820 47346
rect 50428 47292 50820 47294
rect 50428 47282 50484 47292
rect 50764 47282 50820 47292
rect 50316 47068 50484 47124
rect 50428 46676 50484 47068
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50428 46582 50484 46620
rect 50876 46004 50932 48190
rect 51100 47570 51156 47582
rect 51100 47518 51102 47570
rect 51154 47518 51156 47570
rect 48860 43250 48916 43260
rect 49420 43652 49588 43708
rect 49644 45724 49812 45780
rect 50428 45948 50932 46004
rect 50988 47234 51044 47246
rect 50988 47182 50990 47234
rect 51042 47182 51044 47234
rect 48524 43092 48580 43102
rect 47852 42868 47908 42878
rect 47740 42866 47908 42868
rect 47740 42814 47854 42866
rect 47906 42814 47908 42866
rect 47740 42812 47908 42814
rect 47852 42802 47908 42812
rect 47404 42756 47460 42766
rect 47404 41972 47460 42700
rect 47964 41972 48020 41982
rect 47404 41970 47964 41972
rect 47404 41918 47406 41970
rect 47458 41918 47964 41970
rect 47404 41916 47964 41918
rect 47404 41906 47460 41916
rect 47964 41878 48020 41916
rect 48524 41300 48580 43036
rect 49084 41972 49140 41982
rect 48524 41298 48916 41300
rect 48524 41246 48526 41298
rect 48578 41246 48916 41298
rect 48524 41244 48916 41246
rect 48524 41234 48580 41244
rect 48860 41186 48916 41244
rect 48860 41134 48862 41186
rect 48914 41134 48916 41186
rect 48860 41122 48916 41134
rect 47180 40572 47460 40628
rect 46060 39730 46340 39732
rect 46060 39678 46062 39730
rect 46114 39678 46340 39730
rect 46060 39676 46340 39678
rect 46060 39666 46116 39676
rect 45500 38658 45556 38668
rect 46060 37940 46116 37950
rect 45052 37100 45164 37156
rect 44828 36484 44884 36494
rect 44828 36390 44884 36428
rect 44940 36372 44996 36382
rect 45052 36372 45108 37100
rect 45164 37090 45220 37100
rect 45836 37156 45892 37166
rect 45836 37062 45892 37100
rect 45724 36596 45780 36606
rect 45724 36502 45780 36540
rect 44940 36370 45108 36372
rect 44940 36318 44942 36370
rect 44994 36318 45108 36370
rect 44940 36316 45108 36318
rect 45500 36482 45556 36494
rect 45500 36430 45502 36482
rect 45554 36430 45556 36482
rect 44940 36306 44996 36316
rect 45164 36260 45220 36270
rect 45164 36166 45220 36204
rect 44380 33516 44548 33572
rect 44828 35812 44884 35822
rect 44156 32564 44212 32574
rect 44156 32470 44212 32508
rect 44380 31218 44436 33516
rect 44828 33458 44884 35756
rect 45276 35588 45332 35598
rect 45500 35588 45556 36430
rect 45948 36372 46004 36382
rect 45948 36278 46004 36316
rect 45332 35532 45556 35588
rect 45276 35494 45332 35532
rect 45164 35028 45220 35038
rect 45164 34934 45220 34972
rect 45276 34916 45332 34926
rect 45948 34916 46004 34926
rect 45276 34822 45332 34860
rect 45836 34914 46004 34916
rect 45836 34862 45950 34914
rect 46002 34862 46004 34914
rect 45836 34860 46004 34862
rect 46060 34916 46116 37884
rect 46284 37492 46340 39676
rect 46396 39730 46452 39742
rect 46396 39678 46398 39730
rect 46450 39678 46452 39730
rect 46396 39172 46452 39678
rect 46396 39106 46452 39116
rect 47404 38668 47460 40572
rect 48524 40292 48580 40302
rect 48524 39730 48580 40236
rect 48524 39678 48526 39730
rect 48578 39678 48580 39730
rect 48524 39666 48580 39678
rect 49084 39620 49140 41916
rect 49308 41970 49364 41982
rect 49308 41918 49310 41970
rect 49362 41918 49364 41970
rect 49196 41076 49252 41086
rect 49196 40982 49252 41020
rect 49196 39620 49252 39630
rect 49084 39564 49196 39620
rect 49196 39526 49252 39564
rect 49308 39172 49364 41918
rect 47068 38612 47460 38668
rect 48748 39116 49364 39172
rect 46284 37490 46564 37492
rect 46284 37438 46286 37490
rect 46338 37438 46564 37490
rect 46284 37436 46564 37438
rect 46284 37426 46340 37436
rect 46172 37156 46228 37166
rect 46172 36482 46228 37100
rect 46508 36484 46564 37436
rect 46172 36430 46174 36482
rect 46226 36430 46228 36482
rect 46172 36418 46228 36430
rect 46284 36482 46564 36484
rect 46284 36430 46510 36482
rect 46562 36430 46564 36482
rect 46284 36428 46564 36430
rect 46172 35924 46228 35934
rect 46284 35924 46340 36428
rect 46508 36418 46564 36428
rect 46172 35922 46340 35924
rect 46172 35870 46174 35922
rect 46226 35870 46340 35922
rect 46172 35868 46340 35870
rect 46172 35858 46228 35868
rect 46732 35028 46788 35038
rect 46732 34934 46788 34972
rect 46060 34860 46340 34916
rect 45052 34802 45108 34814
rect 45052 34750 45054 34802
rect 45106 34750 45108 34802
rect 45052 34692 45108 34750
rect 45612 34804 45668 34814
rect 45612 34710 45668 34748
rect 45052 33796 45108 34636
rect 45052 33730 45108 33740
rect 44828 33406 44830 33458
rect 44882 33406 44884 33458
rect 44828 33394 44884 33406
rect 44492 33348 44548 33358
rect 44492 32786 44548 33292
rect 45388 33348 45444 33358
rect 45388 33254 45444 33292
rect 44492 32734 44494 32786
rect 44546 32734 44548 32786
rect 44492 32722 44548 32734
rect 45052 33124 45108 33134
rect 45052 32786 45108 33068
rect 45724 33124 45780 33134
rect 45724 33030 45780 33068
rect 45052 32734 45054 32786
rect 45106 32734 45108 32786
rect 45052 32722 45108 32734
rect 44940 32564 44996 32574
rect 44380 31166 44382 31218
rect 44434 31166 44436 31218
rect 44380 31108 44436 31166
rect 44380 31042 44436 31052
rect 44828 31220 44884 31230
rect 44828 31106 44884 31164
rect 44828 31054 44830 31106
rect 44882 31054 44884 31106
rect 44828 31042 44884 31054
rect 44940 30660 44996 32508
rect 45612 32564 45668 32574
rect 45612 32470 45668 32508
rect 45052 32340 45108 32350
rect 45052 32246 45108 32284
rect 45724 31780 45780 31790
rect 45836 31780 45892 34860
rect 45948 34850 46004 34860
rect 46060 33348 46116 33358
rect 46060 33254 46116 33292
rect 45500 31778 45892 31780
rect 45500 31726 45726 31778
rect 45778 31726 45892 31778
rect 45500 31724 45892 31726
rect 45276 31668 45332 31678
rect 45276 31218 45332 31612
rect 45276 31166 45278 31218
rect 45330 31166 45332 31218
rect 45276 31154 45332 31166
rect 45052 31108 45108 31118
rect 45052 31014 45108 31052
rect 45388 30996 45444 31006
rect 44492 30604 44996 30660
rect 45164 30994 45444 30996
rect 45164 30942 45390 30994
rect 45442 30942 45444 30994
rect 45164 30940 45444 30942
rect 44268 27860 44324 27870
rect 44268 27766 44324 27804
rect 44268 26962 44324 26974
rect 44268 26910 44270 26962
rect 44322 26910 44324 26962
rect 44268 26908 44324 26910
rect 44268 26852 44436 26908
rect 44268 26180 44324 26190
rect 44268 26086 44324 26124
rect 44268 25508 44324 25518
rect 44380 25508 44436 26796
rect 44324 25452 44436 25508
rect 44268 25442 44324 25452
rect 44044 25340 44212 25396
rect 43708 24894 43710 24946
rect 43762 24894 43764 24946
rect 43708 24882 43764 24894
rect 43820 24836 43876 24846
rect 43820 24050 43876 24780
rect 43820 23998 43822 24050
rect 43874 23998 43876 24050
rect 43820 23604 43876 23998
rect 43820 23538 43876 23548
rect 44044 24500 44100 24510
rect 43596 23380 43652 23390
rect 44044 23380 44100 24444
rect 43148 23324 43428 23380
rect 43484 23378 43652 23380
rect 43484 23326 43598 23378
rect 43650 23326 43652 23378
rect 43484 23324 43652 23326
rect 43036 23268 43092 23278
rect 43092 23212 43204 23268
rect 43036 23202 43092 23212
rect 43036 23044 43092 23054
rect 43036 22482 43092 22988
rect 43036 22430 43038 22482
rect 43090 22430 43092 22482
rect 43036 22418 43092 22430
rect 42756 21756 42980 21812
rect 42700 21746 42756 21756
rect 42812 21586 42868 21756
rect 42812 21534 42814 21586
rect 42866 21534 42868 21586
rect 42812 21522 42868 21534
rect 43148 21586 43204 23212
rect 43148 21534 43150 21586
rect 43202 21534 43204 21586
rect 42700 21474 42756 21486
rect 42700 21422 42702 21474
rect 42754 21422 42756 21474
rect 42700 21028 42756 21422
rect 43148 21140 43204 21534
rect 43148 21074 43204 21084
rect 42700 20962 42756 20972
rect 43372 20916 43428 23324
rect 43596 23314 43652 23324
rect 43820 23324 44100 23380
rect 43484 23044 43540 23054
rect 43484 22950 43540 22988
rect 43596 22148 43652 22158
rect 43596 22146 43764 22148
rect 43596 22094 43598 22146
rect 43650 22094 43764 22146
rect 43596 22092 43764 22094
rect 43596 22082 43652 22092
rect 43708 22036 43764 22092
rect 43708 21026 43764 21980
rect 43708 20974 43710 21026
rect 43762 20974 43764 21026
rect 43708 20962 43764 20974
rect 43596 20916 43652 20926
rect 43428 20914 43652 20916
rect 43428 20862 43598 20914
rect 43650 20862 43652 20914
rect 43428 20860 43652 20862
rect 43372 20822 43428 20860
rect 43596 20850 43652 20860
rect 42812 20132 42868 20142
rect 42812 20038 42868 20076
rect 43820 20018 43876 23324
rect 43932 23154 43988 23166
rect 43932 23102 43934 23154
rect 43986 23102 43988 23154
rect 43932 21588 43988 23102
rect 44044 23154 44100 23166
rect 44044 23102 44046 23154
rect 44098 23102 44100 23154
rect 44044 22932 44100 23102
rect 44044 22866 44100 22876
rect 44044 22146 44100 22158
rect 44044 22094 44046 22146
rect 44098 22094 44100 22146
rect 44044 22036 44100 22094
rect 44044 21970 44100 21980
rect 44044 21588 44100 21598
rect 43988 21586 44100 21588
rect 43988 21534 44046 21586
rect 44098 21534 44100 21586
rect 43988 21532 44100 21534
rect 43932 21494 43988 21532
rect 44044 21522 44100 21532
rect 43932 21026 43988 21038
rect 43932 20974 43934 21026
rect 43986 20974 43988 21026
rect 43932 20580 43988 20974
rect 44156 20692 44212 25340
rect 44268 25284 44324 25294
rect 44268 24612 44324 25228
rect 44268 24610 44436 24612
rect 44268 24558 44270 24610
rect 44322 24558 44436 24610
rect 44268 24556 44436 24558
rect 44268 24546 44324 24556
rect 44268 23940 44324 23950
rect 44268 23846 44324 23884
rect 44156 20626 44212 20636
rect 44268 23604 44324 23614
rect 43932 20578 44100 20580
rect 43932 20526 43934 20578
rect 43986 20526 44100 20578
rect 43932 20524 44100 20526
rect 43932 20514 43988 20524
rect 44044 20356 44100 20524
rect 44268 20468 44324 23548
rect 44268 20402 44324 20412
rect 44156 20356 44212 20366
rect 44044 20300 44156 20356
rect 44156 20290 44212 20300
rect 43820 19966 43822 20018
rect 43874 19966 43876 20018
rect 42364 19906 42644 19908
rect 42364 19854 42366 19906
rect 42418 19854 42644 19906
rect 42364 19852 42644 19854
rect 43484 19906 43540 19918
rect 43484 19854 43486 19906
rect 43538 19854 43540 19906
rect 42140 19122 42308 19124
rect 42140 19070 42142 19122
rect 42194 19070 42308 19122
rect 42140 19068 42308 19070
rect 42140 19058 42196 19068
rect 41916 18398 41918 18450
rect 41970 18398 41972 18450
rect 41916 18386 41972 18398
rect 42252 17892 42308 19068
rect 42364 19012 42420 19852
rect 43484 19124 43540 19854
rect 43484 19058 43540 19068
rect 43708 19908 43764 19918
rect 42364 18946 42420 18956
rect 42588 18452 42644 18462
rect 42588 18358 42644 18396
rect 43148 18452 43204 18462
rect 43148 18358 43204 18396
rect 43484 18450 43540 18462
rect 43484 18398 43486 18450
rect 43538 18398 43540 18450
rect 42364 18226 42420 18238
rect 42364 18174 42366 18226
rect 42418 18174 42420 18226
rect 42364 18116 42420 18174
rect 43484 18116 43540 18398
rect 42364 18060 43540 18116
rect 42476 17892 42532 17902
rect 42252 17890 42532 17892
rect 42252 17838 42478 17890
rect 42530 17838 42532 17890
rect 42252 17836 42532 17838
rect 42476 17826 42532 17836
rect 43148 17666 43204 18060
rect 43708 17778 43764 19852
rect 43820 19236 43876 19966
rect 43820 19170 43876 19180
rect 43932 20244 43988 20254
rect 43820 19012 43876 19022
rect 43932 19012 43988 20188
rect 44044 20132 44100 20142
rect 44380 20132 44436 24556
rect 44492 21812 44548 30604
rect 45164 30434 45220 30940
rect 45388 30930 45444 30940
rect 45164 30382 45166 30434
rect 45218 30382 45220 30434
rect 45164 30370 45220 30382
rect 45276 30098 45332 30110
rect 45276 30046 45278 30098
rect 45330 30046 45332 30098
rect 45164 29988 45220 29998
rect 45164 29894 45220 29932
rect 44828 29316 44884 29326
rect 44716 29314 44884 29316
rect 44716 29262 44830 29314
rect 44882 29262 44884 29314
rect 44716 29260 44884 29262
rect 44716 28308 44772 29260
rect 44828 29250 44884 29260
rect 44604 27748 44660 27758
rect 44604 27654 44660 27692
rect 44604 26964 44660 26974
rect 44604 26290 44660 26908
rect 44604 26238 44606 26290
rect 44658 26238 44660 26290
rect 44604 26226 44660 26238
rect 44492 21746 44548 21756
rect 44492 21586 44548 21598
rect 44492 21534 44494 21586
rect 44546 21534 44548 21586
rect 44492 21476 44548 21534
rect 44492 20244 44548 21420
rect 44492 20178 44548 20188
rect 44044 20130 44436 20132
rect 44044 20078 44046 20130
rect 44098 20078 44436 20130
rect 44044 20076 44436 20078
rect 44604 20130 44660 20142
rect 44604 20078 44606 20130
rect 44658 20078 44660 20130
rect 44044 19684 44100 20076
rect 44492 20020 44548 20030
rect 44492 19926 44548 19964
rect 44604 19908 44660 20078
rect 44604 19842 44660 19852
rect 44156 19684 44212 19694
rect 44044 19628 44156 19684
rect 44156 19618 44212 19628
rect 44268 19460 44324 19470
rect 43820 19010 43988 19012
rect 43820 18958 43822 19010
rect 43874 18958 43988 19010
rect 43820 18956 43988 18958
rect 43820 18946 43876 18956
rect 43708 17726 43710 17778
rect 43762 17726 43764 17778
rect 43708 17714 43764 17726
rect 43820 18562 43876 18574
rect 43820 18510 43822 18562
rect 43874 18510 43876 18562
rect 43820 18228 43876 18510
rect 43148 17614 43150 17666
rect 43202 17614 43204 17666
rect 43148 17602 43204 17614
rect 42588 17554 42644 17566
rect 43820 17556 43876 18172
rect 42588 17502 42590 17554
rect 42642 17502 42644 17554
rect 41244 17220 41300 17230
rect 41020 16884 41076 16894
rect 41020 15538 41076 16828
rect 41244 16098 41300 17164
rect 42588 17220 42644 17502
rect 43708 17500 43876 17556
rect 42588 17154 42644 17164
rect 42924 17442 42980 17454
rect 42924 17390 42926 17442
rect 42978 17390 42980 17442
rect 42924 17108 42980 17390
rect 42588 16772 42644 16782
rect 42588 16678 42644 16716
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 41244 16034 41300 16046
rect 42028 16210 42084 16222
rect 42028 16158 42030 16210
rect 42082 16158 42084 16210
rect 41020 15486 41022 15538
rect 41074 15486 41076 15538
rect 41020 15474 41076 15486
rect 40908 14578 40964 14588
rect 41356 15202 41412 15214
rect 41356 15150 41358 15202
rect 41410 15150 41412 15202
rect 41356 13860 41412 15150
rect 41916 14420 41972 14430
rect 41916 14326 41972 14364
rect 41356 13794 41412 13804
rect 40908 13636 40964 13646
rect 40908 12962 40964 13580
rect 41804 13636 41860 13646
rect 41804 13542 41860 13580
rect 41804 13412 41860 13422
rect 40908 12910 40910 12962
rect 40962 12910 40964 12962
rect 40908 12898 40964 12910
rect 41020 13074 41076 13086
rect 41020 13022 41022 13074
rect 41074 13022 41076 13074
rect 41020 12964 41076 13022
rect 41020 12898 41076 12908
rect 41020 12738 41076 12750
rect 41020 12686 41022 12738
rect 41074 12686 41076 12738
rect 41020 12068 41076 12686
rect 41020 12002 41076 12012
rect 41468 11396 41524 11406
rect 41580 11396 41636 11406
rect 40796 11394 41300 11396
rect 40796 11342 40798 11394
rect 40850 11342 41300 11394
rect 40796 11340 41300 11342
rect 40796 11330 40852 11340
rect 41020 11172 41076 11182
rect 41020 11078 41076 11116
rect 41020 10948 41076 10958
rect 40460 10836 40516 10846
rect 40460 10742 40516 10780
rect 40908 10164 40964 10174
rect 40908 9714 40964 10108
rect 40908 9662 40910 9714
rect 40962 9662 40964 9714
rect 40908 9650 40964 9662
rect 40796 9604 40852 9614
rect 40684 9602 40852 9604
rect 40684 9550 40798 9602
rect 40850 9550 40852 9602
rect 40684 9548 40852 9550
rect 40684 7364 40740 9548
rect 40796 9538 40852 9548
rect 41020 8932 41076 10892
rect 41132 10610 41188 10622
rect 41132 10558 41134 10610
rect 41186 10558 41188 10610
rect 41132 10052 41188 10558
rect 41132 9986 41188 9996
rect 41244 9828 41300 11340
rect 41468 11394 41580 11396
rect 41468 11342 41470 11394
rect 41522 11342 41580 11394
rect 41468 11340 41580 11342
rect 41468 11330 41524 11340
rect 41356 10836 41412 10846
rect 41356 10742 41412 10780
rect 41468 10612 41524 10622
rect 41468 10518 41524 10556
rect 41580 10164 41636 11340
rect 41692 11170 41748 11182
rect 41692 11118 41694 11170
rect 41746 11118 41748 11170
rect 41692 11060 41748 11118
rect 41692 10994 41748 11004
rect 41804 10276 41860 13356
rect 42028 11396 42084 16158
rect 42364 16100 42420 16110
rect 42364 16006 42420 16044
rect 42700 15428 42756 15438
rect 42476 15204 42532 15214
rect 42252 15092 42532 15148
rect 42252 14754 42308 15092
rect 42252 14702 42254 14754
rect 42306 14702 42308 14754
rect 42252 14690 42308 14702
rect 42700 14644 42756 15372
rect 42364 14642 42756 14644
rect 42364 14590 42702 14642
rect 42754 14590 42756 14642
rect 42364 14588 42756 14590
rect 42252 14532 42308 14542
rect 42364 14532 42420 14588
rect 42700 14578 42756 14588
rect 42252 14530 42420 14532
rect 42252 14478 42254 14530
rect 42306 14478 42420 14530
rect 42252 14476 42420 14478
rect 42252 14466 42308 14476
rect 42588 13636 42644 13646
rect 42588 13186 42644 13580
rect 42588 13134 42590 13186
rect 42642 13134 42644 13186
rect 42588 13122 42644 13134
rect 42476 13076 42532 13086
rect 42252 12964 42308 12974
rect 42252 12870 42308 12908
rect 42476 12850 42532 13020
rect 42476 12798 42478 12850
rect 42530 12798 42532 12850
rect 42476 12786 42532 12798
rect 42028 11330 42084 11340
rect 42700 12068 42756 12078
rect 42028 11170 42084 11182
rect 42028 11118 42030 11170
rect 42082 11118 42084 11170
rect 41916 11060 41972 11070
rect 41916 10834 41972 11004
rect 41916 10782 41918 10834
rect 41970 10782 41972 10834
rect 41916 10770 41972 10782
rect 42028 10724 42084 11118
rect 42028 10658 42084 10668
rect 42140 11172 42196 11182
rect 42140 10722 42196 11116
rect 42140 10670 42142 10722
rect 42194 10670 42196 10722
rect 42140 10612 42196 10670
rect 42364 11170 42420 11182
rect 42364 11118 42366 11170
rect 42418 11118 42420 11170
rect 42252 10612 42308 10622
rect 42140 10556 42252 10612
rect 42252 10546 42308 10556
rect 41916 10500 41972 10510
rect 41972 10444 42084 10500
rect 41916 10406 41972 10444
rect 41804 10220 41972 10276
rect 41580 10108 41860 10164
rect 41356 9828 41412 9838
rect 41244 9826 41412 9828
rect 41244 9774 41358 9826
rect 41410 9774 41412 9826
rect 41244 9772 41412 9774
rect 41356 9762 41412 9772
rect 41804 9826 41860 10108
rect 41804 9774 41806 9826
rect 41858 9774 41860 9826
rect 41804 9762 41860 9774
rect 41020 8876 41524 8932
rect 41468 8258 41524 8876
rect 41468 8206 41470 8258
rect 41522 8206 41524 8258
rect 40684 7298 40740 7308
rect 40796 8036 40852 8046
rect 40796 6690 40852 7980
rect 41244 7924 41300 7934
rect 40796 6638 40798 6690
rect 40850 6638 40852 6690
rect 40796 6626 40852 6638
rect 40908 7698 40964 7710
rect 40908 7646 40910 7698
rect 40962 7646 40964 7698
rect 40908 6578 40964 7646
rect 41244 7474 41300 7868
rect 41468 7700 41524 8206
rect 41468 7634 41524 7644
rect 41804 8148 41860 8158
rect 41916 8148 41972 10220
rect 42028 9268 42084 10444
rect 42364 10164 42420 11118
rect 42700 10500 42756 12012
rect 42924 11844 42980 17052
rect 43148 17444 43204 17454
rect 43148 16882 43204 17388
rect 43148 16830 43150 16882
rect 43202 16830 43204 16882
rect 43148 16818 43204 16830
rect 43484 15204 43540 15242
rect 43484 15138 43540 15148
rect 43036 13076 43092 13086
rect 43036 12982 43092 13020
rect 42924 11778 42980 11788
rect 42812 11172 42868 11182
rect 43260 11172 43316 11182
rect 42812 11170 43316 11172
rect 42812 11118 42814 11170
rect 42866 11118 43262 11170
rect 43314 11118 43316 11170
rect 42812 11116 43316 11118
rect 42812 10724 42868 11116
rect 43260 11106 43316 11116
rect 43372 11060 43428 11070
rect 42868 10668 42980 10724
rect 42812 10658 42868 10668
rect 42924 10610 42980 10668
rect 42924 10558 42926 10610
rect 42978 10558 42980 10610
rect 42924 10546 42980 10558
rect 43372 10610 43428 11004
rect 43708 10836 43764 17500
rect 43932 17220 43988 18956
rect 43820 16324 43876 16334
rect 43820 16098 43876 16268
rect 43820 16046 43822 16098
rect 43874 16046 43876 16098
rect 43820 16034 43876 16046
rect 43932 14420 43988 17164
rect 43932 14354 43988 14364
rect 44044 19404 44268 19460
rect 43932 13636 43988 13646
rect 43932 13542 43988 13580
rect 43708 10770 43764 10780
rect 43372 10558 43374 10610
rect 43426 10558 43428 10610
rect 43372 10546 43428 10558
rect 43820 10612 43876 10622
rect 43820 10518 43876 10556
rect 42700 10444 42868 10500
rect 42364 10098 42420 10108
rect 42700 9604 42756 9614
rect 42252 9268 42308 9278
rect 42028 9266 42308 9268
rect 42028 9214 42254 9266
rect 42306 9214 42308 9266
rect 42028 9212 42308 9214
rect 42252 9202 42308 9212
rect 42140 9042 42196 9054
rect 42140 8990 42142 9042
rect 42194 8990 42196 9042
rect 42140 8484 42196 8990
rect 42476 9044 42532 9054
rect 42476 8950 42532 8988
rect 42140 8418 42196 8428
rect 42700 8258 42756 9548
rect 42812 8930 42868 10444
rect 43932 10386 43988 10398
rect 43932 10334 43934 10386
rect 43986 10334 43988 10386
rect 43932 9828 43988 10334
rect 43596 9714 43652 9726
rect 43596 9662 43598 9714
rect 43650 9662 43652 9714
rect 43596 9604 43652 9662
rect 43596 9538 43652 9548
rect 42812 8878 42814 8930
rect 42866 8878 42868 8930
rect 42812 8484 42868 8878
rect 42812 8418 42868 8428
rect 43820 9268 43876 9278
rect 43148 8372 43204 8382
rect 42700 8206 42702 8258
rect 42754 8206 42756 8258
rect 42700 8194 42756 8206
rect 42924 8260 42980 8270
rect 42924 8166 42980 8204
rect 43148 8258 43204 8316
rect 43148 8206 43150 8258
rect 43202 8206 43204 8258
rect 43148 8194 43204 8206
rect 43820 8260 43876 9212
rect 43820 8194 43876 8204
rect 43932 8258 43988 9772
rect 43932 8206 43934 8258
rect 43986 8206 43988 8258
rect 43932 8194 43988 8206
rect 44044 8372 44100 19404
rect 44268 19394 44324 19404
rect 44268 19012 44324 19022
rect 44156 17556 44212 17566
rect 44156 17462 44212 17500
rect 44156 16772 44212 16782
rect 44156 15316 44212 16716
rect 44268 16660 44324 18956
rect 44492 18340 44548 18350
rect 44492 16882 44548 18284
rect 44604 18338 44660 18350
rect 44604 18286 44606 18338
rect 44658 18286 44660 18338
rect 44604 17332 44660 18286
rect 44604 17266 44660 17276
rect 44492 16830 44494 16882
rect 44546 16830 44548 16882
rect 44492 16818 44548 16830
rect 44268 16594 44324 16604
rect 44716 16324 44772 28252
rect 45276 28084 45332 30046
rect 45500 29652 45556 31724
rect 45724 31714 45780 31724
rect 45724 29988 45780 29998
rect 45724 29894 45780 29932
rect 45500 29558 45556 29596
rect 45388 28084 45444 28094
rect 45276 28082 45444 28084
rect 45276 28030 45390 28082
rect 45442 28030 45444 28082
rect 45276 28028 45444 28030
rect 45388 28018 45444 28028
rect 45612 27970 45668 27982
rect 45612 27918 45614 27970
rect 45666 27918 45668 27970
rect 45052 27860 45108 27870
rect 45108 27804 45332 27860
rect 45052 27766 45108 27804
rect 45052 27300 45108 27310
rect 45052 27206 45108 27244
rect 44828 27074 44884 27086
rect 44828 27022 44830 27074
rect 44882 27022 44884 27074
rect 44828 26852 44884 27022
rect 44828 26786 44884 26796
rect 45164 26404 45220 26414
rect 45164 26310 45220 26348
rect 44828 24610 44884 24622
rect 44828 24558 44830 24610
rect 44882 24558 44884 24610
rect 44828 24500 44884 24558
rect 44828 24434 44884 24444
rect 44940 24052 44996 24062
rect 45276 24052 45332 27804
rect 45612 27524 45668 27918
rect 45612 27458 45668 27468
rect 45724 27858 45780 27870
rect 45724 27806 45726 27858
rect 45778 27806 45780 27858
rect 45388 27300 45444 27310
rect 45724 27300 45780 27806
rect 45388 27298 45780 27300
rect 45388 27246 45390 27298
rect 45442 27246 45726 27298
rect 45778 27246 45780 27298
rect 45388 27244 45780 27246
rect 45388 27234 45444 27244
rect 45724 27206 45780 27244
rect 45948 27524 46004 27534
rect 45948 27186 46004 27468
rect 45948 27134 45950 27186
rect 46002 27134 46004 27186
rect 45948 27122 46004 27134
rect 44940 24050 45332 24052
rect 44940 23998 44942 24050
rect 44994 23998 45332 24050
rect 44940 23996 45332 23998
rect 44940 23986 44996 23996
rect 45052 23940 45108 23996
rect 44940 23380 44996 23390
rect 44828 23324 44940 23380
rect 44828 22370 44884 23324
rect 44940 23314 44996 23324
rect 44940 23156 44996 23166
rect 45052 23156 45108 23884
rect 45276 23938 45332 23996
rect 45276 23886 45278 23938
rect 45330 23886 45332 23938
rect 45276 23874 45332 23886
rect 45388 26180 45444 26190
rect 45388 24722 45444 26124
rect 46284 24836 46340 34860
rect 46396 31668 46452 31678
rect 46396 31574 46452 31612
rect 46508 29428 46564 29438
rect 46844 29428 46900 29438
rect 47068 29428 47124 38612
rect 48188 37268 48244 37278
rect 48188 37174 48244 37212
rect 47292 36596 47348 36606
rect 47292 36502 47348 36540
rect 47180 36260 47236 36270
rect 47180 33572 47236 36204
rect 48748 34356 48804 39116
rect 49420 39060 49476 43652
rect 49644 40404 49700 45724
rect 50316 45106 50372 45118
rect 50316 45054 50318 45106
rect 50370 45054 50372 45106
rect 49980 44996 50036 45006
rect 50316 44996 50372 45054
rect 49980 44994 50372 44996
rect 49980 44942 49982 44994
rect 50034 44942 50372 44994
rect 49980 44940 50372 44942
rect 49980 44930 50036 44940
rect 49756 44100 49812 44110
rect 49756 42194 49812 44044
rect 49868 43316 49924 43326
rect 49924 43260 50036 43316
rect 49868 43250 49924 43260
rect 49980 42866 50036 43260
rect 49980 42814 49982 42866
rect 50034 42814 50036 42866
rect 49980 42802 50036 42814
rect 49756 42142 49758 42194
rect 49810 42142 49812 42194
rect 49756 40516 49812 42142
rect 49868 42644 49924 42654
rect 49868 41970 49924 42588
rect 49980 42084 50036 42094
rect 49980 41990 50036 42028
rect 49868 41918 49870 41970
rect 49922 41918 49924 41970
rect 49868 41906 49924 41918
rect 50316 41972 50372 44940
rect 50428 42084 50484 45948
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50876 44098 50932 44110
rect 50876 44046 50878 44098
rect 50930 44046 50932 44098
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50876 43764 50932 44046
rect 50876 43698 50932 43708
rect 50988 43876 51044 47182
rect 51100 46786 51156 47518
rect 51100 46734 51102 46786
rect 51154 46734 51156 46786
rect 51100 46722 51156 46734
rect 51100 44996 51156 45006
rect 51996 44996 52052 50542
rect 53228 49924 53284 49934
rect 53228 49698 53284 49868
rect 53228 49646 53230 49698
rect 53282 49646 53284 49698
rect 53228 49634 53284 49646
rect 53004 48018 53060 48030
rect 53004 47966 53006 48018
rect 53058 47966 53060 48018
rect 53004 46228 53060 47966
rect 53228 46564 53284 46574
rect 53228 46470 53284 46508
rect 53004 46162 53060 46172
rect 51100 44994 51828 44996
rect 51100 44942 51102 44994
rect 51154 44942 51828 44994
rect 51100 44940 51828 44942
rect 51100 44930 51156 44940
rect 51100 44772 51156 44782
rect 51100 44322 51156 44716
rect 51772 44434 51828 44940
rect 51996 44930 52052 44940
rect 53228 44996 53284 45006
rect 53228 44902 53284 44940
rect 51772 44382 51774 44434
rect 51826 44382 51828 44434
rect 51772 44370 51828 44382
rect 51100 44270 51102 44322
rect 51154 44270 51156 44322
rect 51100 44258 51156 44270
rect 51212 44324 51268 44334
rect 51660 44324 51716 44334
rect 51212 44322 51716 44324
rect 51212 44270 51214 44322
rect 51266 44270 51662 44322
rect 51714 44270 51716 44322
rect 51212 44268 51716 44270
rect 51212 44258 51268 44268
rect 51660 44258 51716 44268
rect 51324 44100 51380 44110
rect 51324 44006 51380 44044
rect 51884 44098 51940 44110
rect 51884 44046 51886 44098
rect 51938 44046 51940 44098
rect 51884 43876 51940 44046
rect 50988 43820 51940 43876
rect 50988 43092 51044 43820
rect 51100 43540 51156 43550
rect 53004 43540 53060 43550
rect 51100 43538 51268 43540
rect 51100 43486 51102 43538
rect 51154 43486 51268 43538
rect 51100 43484 51268 43486
rect 51100 43474 51156 43484
rect 50876 43036 51044 43092
rect 50652 42644 50708 42654
rect 50652 42550 50708 42588
rect 50876 42642 50932 43036
rect 50876 42590 50878 42642
rect 50930 42590 50932 42642
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50428 42018 50484 42028
rect 50316 41878 50372 41916
rect 49980 41188 50036 41198
rect 49980 41186 50260 41188
rect 49980 41134 49982 41186
rect 50034 41134 50260 41186
rect 49980 41132 50260 41134
rect 49980 41122 50036 41132
rect 49756 40460 50148 40516
rect 49644 40348 50036 40404
rect 49868 39508 49924 39518
rect 49196 39004 49476 39060
rect 49644 39396 49700 39406
rect 49196 38668 49252 39004
rect 48972 38612 49252 38668
rect 49308 38834 49364 38846
rect 49308 38782 49310 38834
rect 49362 38782 49364 38834
rect 48972 37268 49028 38612
rect 49308 37716 49364 38782
rect 49308 37650 49364 37660
rect 49420 38052 49476 38062
rect 49420 37492 49476 37996
rect 48860 35364 48916 35374
rect 48860 35026 48916 35308
rect 48860 34974 48862 35026
rect 48914 34974 48916 35026
rect 48860 34962 48916 34974
rect 48748 34290 48804 34300
rect 48860 34020 48916 34030
rect 48972 34020 49028 37212
rect 49308 37490 49476 37492
rect 49308 37438 49422 37490
rect 49474 37438 49476 37490
rect 49308 37436 49476 37438
rect 49196 35588 49252 35598
rect 49196 35494 49252 35532
rect 49308 34916 49364 37436
rect 49420 37426 49476 37436
rect 49644 37490 49700 39340
rect 49868 39058 49924 39452
rect 49868 39006 49870 39058
rect 49922 39006 49924 39058
rect 49868 38994 49924 39006
rect 49980 39060 50036 40348
rect 49980 38966 50036 39004
rect 49756 38834 49812 38846
rect 49756 38782 49758 38834
rect 49810 38782 49812 38834
rect 49756 38052 49812 38782
rect 49756 37986 49812 37996
rect 49980 38836 50036 38846
rect 49980 38162 50036 38780
rect 49980 38110 49982 38162
rect 50034 38110 50036 38162
rect 49644 37438 49646 37490
rect 49698 37438 49700 37490
rect 49532 37156 49588 37166
rect 49532 37062 49588 37100
rect 49420 36596 49476 36606
rect 49644 36596 49700 37438
rect 49420 36594 49700 36596
rect 49420 36542 49422 36594
rect 49474 36542 49700 36594
rect 49420 36540 49700 36542
rect 49420 36530 49476 36540
rect 49756 36372 49812 36382
rect 49756 35364 49812 36316
rect 49980 35924 50036 38110
rect 49980 35830 50036 35868
rect 50092 36484 50148 40460
rect 49532 34916 49588 34926
rect 48636 33964 48860 34020
rect 48916 33964 49028 34020
rect 49084 34914 49588 34916
rect 49084 34862 49534 34914
rect 49586 34862 49588 34914
rect 49084 34860 49588 34862
rect 47180 33506 47236 33516
rect 47292 33796 47348 33806
rect 46508 29426 47068 29428
rect 46508 29374 46510 29426
rect 46562 29374 46846 29426
rect 46898 29374 47068 29426
rect 46508 29372 47068 29374
rect 46508 29362 46564 29372
rect 46844 29362 46900 29372
rect 47068 29362 47124 29372
rect 47292 29316 47348 33740
rect 48524 31890 48580 31902
rect 48524 31838 48526 31890
rect 48578 31838 48580 31890
rect 48300 29988 48356 29998
rect 48524 29988 48580 31838
rect 48356 29932 48580 29988
rect 47404 29540 47460 29550
rect 47852 29540 47908 29550
rect 47404 29538 47908 29540
rect 47404 29486 47406 29538
rect 47458 29486 47854 29538
rect 47906 29486 47908 29538
rect 47404 29484 47908 29486
rect 47404 29474 47460 29484
rect 47852 29474 47908 29484
rect 48188 29540 48244 29550
rect 48188 29446 48244 29484
rect 47964 29428 48020 29438
rect 48020 29372 48132 29428
rect 47292 29260 47460 29316
rect 47068 29202 47124 29214
rect 47068 29150 47070 29202
rect 47122 29150 47124 29202
rect 47068 29092 47124 29150
rect 47404 29204 47460 29260
rect 47964 29204 48020 29372
rect 48076 29316 48132 29372
rect 48076 29260 48244 29316
rect 47404 29148 47572 29204
rect 47068 29036 47460 29092
rect 47068 28868 47124 28878
rect 47068 28774 47124 28812
rect 47404 28866 47460 29036
rect 47404 28814 47406 28866
rect 47458 28814 47460 28866
rect 47404 28802 47460 28814
rect 47516 28644 47572 29148
rect 47292 28588 47572 28644
rect 47628 29148 48020 29204
rect 46508 28532 46564 28542
rect 46508 28438 46564 28476
rect 46732 28530 46788 28542
rect 46732 28478 46734 28530
rect 46786 28478 46788 28530
rect 46732 28082 46788 28478
rect 46732 28030 46734 28082
rect 46786 28030 46788 28082
rect 46732 28018 46788 28030
rect 46508 27972 46564 27982
rect 46508 27970 46676 27972
rect 46508 27918 46510 27970
rect 46562 27918 46676 27970
rect 46508 27916 46676 27918
rect 46508 27906 46564 27916
rect 46396 27858 46452 27870
rect 46396 27806 46398 27858
rect 46450 27806 46452 27858
rect 46396 27298 46452 27806
rect 46396 27246 46398 27298
rect 46450 27246 46452 27298
rect 46396 27234 46452 27246
rect 46620 27300 46676 27916
rect 47068 27300 47124 27310
rect 46620 27244 47068 27300
rect 46508 27188 46564 27198
rect 46564 27132 46676 27188
rect 46508 27122 46564 27132
rect 46620 27074 46676 27132
rect 46620 27022 46622 27074
rect 46674 27022 46676 27074
rect 46620 26908 46676 27022
rect 47068 27074 47124 27244
rect 47068 27022 47070 27074
rect 47122 27022 47124 27074
rect 47068 27010 47124 27022
rect 47292 26908 47348 28588
rect 47628 28084 47684 29148
rect 47964 28868 48020 28878
rect 47964 28642 48020 28812
rect 47964 28590 47966 28642
rect 48018 28590 48020 28642
rect 47964 28578 48020 28590
rect 48188 28642 48244 29260
rect 48188 28590 48190 28642
rect 48242 28590 48244 28642
rect 48188 28578 48244 28590
rect 48300 28756 48356 29932
rect 48300 28642 48356 28700
rect 48300 28590 48302 28642
rect 48354 28590 48356 28642
rect 48300 28578 48356 28590
rect 46620 26852 46900 26908
rect 46284 24770 46340 24780
rect 45388 24670 45390 24722
rect 45442 24670 45444 24722
rect 45388 23380 45444 24670
rect 46060 24612 46116 24622
rect 46060 24610 46676 24612
rect 46060 24558 46062 24610
rect 46114 24558 46676 24610
rect 46060 24556 46676 24558
rect 46060 24546 46116 24556
rect 46620 24162 46676 24556
rect 46620 24110 46622 24162
rect 46674 24110 46676 24162
rect 46620 24098 46676 24110
rect 46284 23828 46340 23838
rect 46172 23772 46284 23828
rect 45612 23716 45668 23726
rect 45724 23716 45780 23726
rect 45612 23714 45724 23716
rect 45612 23662 45614 23714
rect 45666 23662 45724 23714
rect 45612 23660 45724 23662
rect 45612 23650 45668 23660
rect 45388 23314 45444 23324
rect 44940 23154 45108 23156
rect 44940 23102 44942 23154
rect 44994 23102 45108 23154
rect 44940 23100 45108 23102
rect 44940 23090 44996 23100
rect 45388 23042 45444 23054
rect 45388 22990 45390 23042
rect 45442 22990 45444 23042
rect 45388 22932 45444 22990
rect 45388 22866 45444 22876
rect 44828 22318 44830 22370
rect 44882 22318 44884 22370
rect 44828 22306 44884 22318
rect 45612 22258 45668 22270
rect 45612 22206 45614 22258
rect 45666 22206 45668 22258
rect 45052 21476 45108 21486
rect 45052 21382 45108 21420
rect 44940 20802 44996 20814
rect 44940 20750 44942 20802
rect 44994 20750 44996 20802
rect 44940 20356 44996 20750
rect 45164 20804 45220 20814
rect 45164 20710 45220 20748
rect 45388 20804 45444 20814
rect 45388 20710 45444 20748
rect 45052 20580 45108 20590
rect 45612 20580 45668 22206
rect 45052 20578 45668 20580
rect 45052 20526 45054 20578
rect 45106 20526 45668 20578
rect 45052 20524 45668 20526
rect 45052 20514 45108 20524
rect 44940 20290 44996 20300
rect 45500 20356 45556 20366
rect 45388 20244 45444 20254
rect 44828 20130 44884 20142
rect 44828 20078 44830 20130
rect 44882 20078 44884 20130
rect 44828 20020 44884 20078
rect 45052 20132 45108 20142
rect 44940 20020 44996 20030
rect 44828 20018 44996 20020
rect 44828 19966 44942 20018
rect 44994 19966 44996 20018
rect 44828 19964 44996 19966
rect 44940 19954 44996 19964
rect 44940 19684 44996 19694
rect 44940 19010 44996 19628
rect 44940 18958 44942 19010
rect 44994 18958 44996 19010
rect 44940 18676 44996 18958
rect 44716 16230 44772 16268
rect 44828 18620 44996 18676
rect 44268 16212 44324 16222
rect 44268 16118 44324 16156
rect 44716 15316 44772 15326
rect 44156 15314 44772 15316
rect 44156 15262 44158 15314
rect 44210 15262 44718 15314
rect 44770 15262 44772 15314
rect 44156 15260 44772 15262
rect 44156 15250 44212 15260
rect 41804 8146 41972 8148
rect 41804 8094 41806 8146
rect 41858 8094 41972 8146
rect 41804 8092 41972 8094
rect 43372 8146 43428 8158
rect 43372 8094 43374 8146
rect 43426 8094 43428 8146
rect 41244 7422 41246 7474
rect 41298 7422 41300 7474
rect 41244 7410 41300 7422
rect 41692 7476 41748 7486
rect 41804 7476 41860 8092
rect 42588 8036 42644 8046
rect 42588 7942 42644 7980
rect 43372 8036 43428 8094
rect 43708 8036 43764 8046
rect 44044 8036 44100 8316
rect 43372 8034 43764 8036
rect 43372 7982 43710 8034
rect 43762 7982 43764 8034
rect 43372 7980 43764 7982
rect 42140 7700 42196 7710
rect 42140 7606 42196 7644
rect 41692 7474 41860 7476
rect 41692 7422 41694 7474
rect 41746 7422 41860 7474
rect 41692 7420 41860 7422
rect 42476 7586 42532 7598
rect 42476 7534 42478 7586
rect 42530 7534 42532 7586
rect 41692 7410 41748 7420
rect 41020 7252 41076 7262
rect 41020 7158 41076 7196
rect 41804 7252 41860 7262
rect 41804 6804 41860 7196
rect 42476 6916 42532 7534
rect 43036 7362 43092 7374
rect 43036 7310 43038 7362
rect 43090 7310 43092 7362
rect 43036 7252 43092 7310
rect 43036 7186 43092 7196
rect 42476 6850 42532 6860
rect 43372 6804 43428 7980
rect 43708 7970 43764 7980
rect 43820 7980 44100 8036
rect 44156 14980 44212 14990
rect 43708 7700 43764 7710
rect 43820 7700 43876 7980
rect 43708 7698 43876 7700
rect 43708 7646 43710 7698
rect 43762 7646 43876 7698
rect 43708 7644 43876 7646
rect 43708 7634 43764 7644
rect 43820 6916 43876 6926
rect 43820 6822 43876 6860
rect 41804 6748 42084 6804
rect 40908 6526 40910 6578
rect 40962 6526 40964 6578
rect 40908 6514 40964 6526
rect 41132 6468 41188 6478
rect 41132 6466 41972 6468
rect 41132 6414 41134 6466
rect 41186 6414 41972 6466
rect 41132 6412 41972 6414
rect 41132 6402 41188 6412
rect 40908 5236 40964 5246
rect 40908 5142 40964 5180
rect 41356 4898 41412 4910
rect 41356 4846 41358 4898
rect 41410 4846 41412 4898
rect 41244 4340 41300 4350
rect 41356 4340 41412 4846
rect 41916 4450 41972 6412
rect 41916 4398 41918 4450
rect 41970 4398 41972 4450
rect 41916 4386 41972 4398
rect 41300 4284 41412 4340
rect 41244 4246 41300 4284
rect 40236 3614 40238 3666
rect 40290 3614 40292 3666
rect 40236 3602 40292 3614
rect 41356 3668 41412 4284
rect 42028 4228 42084 6748
rect 43372 6690 43428 6748
rect 43372 6638 43374 6690
rect 43426 6638 43428 6690
rect 43372 6626 43428 6638
rect 43596 6692 43652 6702
rect 43596 6598 43652 6636
rect 44044 6690 44100 6702
rect 44044 6638 44046 6690
rect 44098 6638 44100 6690
rect 44044 6468 44100 6638
rect 44044 6402 44100 6412
rect 42028 4162 42084 4172
rect 43708 4564 43764 4574
rect 41356 3602 41412 3612
rect 42028 3668 42084 3678
rect 42028 3574 42084 3612
rect 43708 3668 43764 4508
rect 44044 4228 44100 4238
rect 44044 4134 44100 4172
rect 35532 3556 35588 3566
rect 35532 3462 35588 3500
rect 35980 3556 36036 3566
rect 35980 3462 36036 3500
rect 43708 3554 43764 3612
rect 43708 3502 43710 3554
rect 43762 3502 43764 3554
rect 43708 3490 43764 3502
rect 38556 3444 38612 3454
rect 38556 800 38612 3388
rect 39340 3444 39396 3482
rect 39340 3378 39396 3388
rect 39788 3444 39844 3482
rect 39788 3378 39844 3388
rect 42476 3444 42532 3454
rect 42700 3444 42756 3454
rect 42476 3442 42756 3444
rect 42476 3390 42478 3442
rect 42530 3390 42702 3442
rect 42754 3390 42756 3442
rect 42476 3388 42756 3390
rect 43036 3444 43092 3482
rect 42476 3378 42532 3388
rect 42700 3332 42868 3388
rect 43036 3378 43092 3388
rect 44156 3444 44212 14924
rect 44604 14644 44660 15260
rect 44716 15250 44772 15260
rect 44716 14980 44772 14990
rect 44828 14980 44884 18620
rect 45052 17556 45108 20076
rect 45388 20130 45444 20188
rect 45388 20078 45390 20130
rect 45442 20078 45444 20130
rect 45388 20066 45444 20078
rect 45500 20130 45556 20300
rect 45500 20078 45502 20130
rect 45554 20078 45556 20130
rect 45500 20066 45556 20078
rect 45612 20020 45668 20030
rect 45388 19012 45444 19022
rect 45388 18918 45444 18956
rect 45612 18788 45668 19964
rect 45388 18732 45668 18788
rect 45164 18450 45220 18462
rect 45164 18398 45166 18450
rect 45218 18398 45220 18450
rect 45164 17780 45220 18398
rect 45164 17714 45220 17724
rect 45052 17500 45220 17556
rect 44940 17442 44996 17454
rect 44940 17390 44942 17442
rect 44994 17390 44996 17442
rect 44940 17220 44996 17390
rect 44940 17154 44996 17164
rect 45052 16996 45108 17006
rect 45052 16902 45108 16940
rect 44940 16322 44996 16334
rect 44940 16270 44942 16322
rect 44994 16270 44996 16322
rect 44940 16210 44996 16270
rect 44940 16158 44942 16210
rect 44994 16158 44996 16210
rect 44940 16146 44996 16158
rect 44772 14924 44884 14980
rect 44716 14914 44772 14924
rect 44604 14588 44772 14644
rect 44716 13748 44772 14588
rect 45164 13972 45220 17500
rect 45276 15316 45332 15326
rect 45276 14532 45332 15260
rect 45388 14756 45444 18732
rect 45500 17556 45556 17566
rect 45500 17442 45556 17500
rect 45500 17390 45502 17442
rect 45554 17390 45556 17442
rect 45500 16884 45556 17390
rect 45500 16818 45556 16828
rect 45724 16548 45780 23660
rect 45948 20804 46004 20814
rect 45836 19348 45892 19358
rect 45948 19348 46004 20748
rect 46060 19908 46116 19918
rect 46060 19814 46116 19852
rect 45892 19292 46004 19348
rect 45836 19282 45892 19292
rect 45948 17668 46004 17678
rect 45948 17574 46004 17612
rect 45724 16492 46116 16548
rect 45500 15540 45556 15550
rect 45500 15446 45556 15484
rect 45836 15316 45892 15354
rect 45836 15250 45892 15260
rect 45388 14690 45444 14700
rect 45948 14756 46004 14766
rect 45836 14644 45892 14654
rect 45388 14532 45444 14542
rect 45276 14530 45444 14532
rect 45276 14478 45390 14530
rect 45442 14478 45444 14530
rect 45276 14476 45444 14478
rect 45164 13916 45332 13972
rect 45164 13748 45220 13758
rect 44716 13746 45220 13748
rect 44716 13694 44718 13746
rect 44770 13694 45166 13746
rect 45218 13694 45220 13746
rect 44716 13692 45220 13694
rect 44604 13524 44660 13534
rect 44604 12402 44660 13468
rect 44604 12350 44606 12402
rect 44658 12350 44660 12402
rect 44604 12338 44660 12350
rect 44268 6580 44324 6590
rect 44268 6486 44324 6524
rect 44380 6466 44436 6478
rect 44380 6414 44382 6466
rect 44434 6414 44436 6466
rect 44380 5236 44436 6414
rect 44716 5684 44772 13692
rect 45164 13682 45220 13692
rect 44940 12404 44996 12414
rect 44940 12402 45220 12404
rect 44940 12350 44942 12402
rect 44994 12350 45220 12402
rect 44940 12348 45220 12350
rect 44940 12338 44996 12348
rect 44828 12178 44884 12190
rect 44828 12126 44830 12178
rect 44882 12126 44884 12178
rect 44828 11060 44884 12126
rect 45052 12178 45108 12190
rect 45052 12126 45054 12178
rect 45106 12126 45108 12178
rect 44828 10994 44884 11004
rect 44940 11172 44996 11182
rect 44940 10050 44996 11116
rect 45052 10612 45108 12126
rect 45164 11394 45220 12348
rect 45164 11342 45166 11394
rect 45218 11342 45220 11394
rect 45164 11330 45220 11342
rect 45052 10498 45108 10556
rect 45164 11060 45220 11070
rect 45164 10610 45220 11004
rect 45164 10558 45166 10610
rect 45218 10558 45220 10610
rect 45164 10546 45220 10558
rect 45052 10446 45054 10498
rect 45106 10446 45108 10498
rect 45052 10434 45108 10446
rect 45276 10052 45332 13916
rect 45388 13412 45444 14476
rect 45388 13346 45444 13356
rect 45836 13076 45892 14588
rect 45948 13524 46004 14700
rect 45948 13458 46004 13468
rect 45836 13010 45892 13020
rect 46060 12402 46116 16492
rect 46172 15540 46228 23772
rect 46284 23734 46340 23772
rect 46732 23828 46788 23838
rect 46732 23734 46788 23772
rect 46732 21700 46788 21710
rect 46284 20692 46340 20702
rect 46284 20018 46340 20636
rect 46732 20244 46788 21644
rect 46732 20130 46788 20188
rect 46732 20078 46734 20130
rect 46786 20078 46788 20130
rect 46732 20066 46788 20078
rect 46844 20132 46900 26852
rect 47180 26852 47348 26908
rect 47404 28082 47684 28084
rect 47404 28030 47630 28082
rect 47682 28030 47684 28082
rect 47404 28028 47684 28030
rect 46956 25284 47012 25294
rect 46956 24162 47012 25228
rect 46956 24110 46958 24162
rect 47010 24110 47012 24162
rect 46956 24098 47012 24110
rect 47180 22148 47236 26852
rect 47404 23716 47460 28028
rect 47628 28018 47684 28028
rect 48076 28532 48132 28542
rect 48076 28084 48132 28476
rect 48076 28082 48580 28084
rect 48076 28030 48078 28082
rect 48130 28030 48580 28082
rect 48076 28028 48580 28030
rect 48076 28018 48132 28028
rect 48412 27748 48468 27758
rect 47628 27524 47684 27534
rect 47516 27300 47572 27310
rect 47516 27206 47572 27244
rect 47628 27186 47684 27468
rect 47628 27134 47630 27186
rect 47682 27134 47684 27186
rect 47628 26908 47684 27134
rect 47404 23650 47460 23660
rect 47516 26852 48132 26908
rect 47180 22082 47236 22092
rect 47516 21028 47572 26852
rect 48076 26850 48132 26852
rect 48076 26798 48078 26850
rect 48130 26798 48132 26850
rect 48076 26786 48132 26798
rect 48412 25282 48468 27692
rect 48412 25230 48414 25282
rect 48466 25230 48468 25282
rect 48188 24612 48244 24622
rect 48188 23716 48244 24556
rect 48188 23714 48356 23716
rect 48188 23662 48190 23714
rect 48242 23662 48356 23714
rect 48188 23660 48356 23662
rect 48188 23650 48244 23660
rect 47964 23042 48020 23054
rect 47964 22990 47966 23042
rect 48018 22990 48020 23042
rect 47740 22482 47796 22494
rect 47740 22430 47742 22482
rect 47794 22430 47796 22482
rect 47740 21700 47796 22430
rect 47964 22484 48020 22990
rect 47964 22418 48020 22428
rect 47740 21634 47796 21644
rect 48076 22370 48132 22382
rect 48076 22318 48078 22370
rect 48130 22318 48132 22370
rect 47740 21476 47796 21486
rect 48076 21476 48132 22318
rect 47740 21474 48132 21476
rect 47740 21422 47742 21474
rect 47794 21422 48132 21474
rect 47740 21420 48132 21422
rect 47516 20972 47684 21028
rect 47404 20244 47460 20254
rect 46284 19966 46286 20018
rect 46338 19966 46340 20018
rect 46284 18340 46340 19966
rect 46508 19906 46564 19918
rect 46508 19854 46510 19906
rect 46562 19854 46564 19906
rect 46508 18564 46564 19854
rect 46844 19348 46900 20076
rect 46956 20242 47460 20244
rect 46956 20190 47406 20242
rect 47458 20190 47460 20242
rect 46956 20188 47460 20190
rect 46956 20130 47012 20188
rect 47404 20178 47460 20188
rect 46956 20078 46958 20130
rect 47010 20078 47012 20130
rect 46956 20066 47012 20078
rect 47516 20132 47572 20142
rect 47516 20038 47572 20076
rect 47292 20020 47348 20030
rect 47292 19926 47348 19964
rect 47068 19348 47124 19358
rect 46844 19346 47124 19348
rect 46844 19294 47070 19346
rect 47122 19294 47124 19346
rect 46844 19292 47124 19294
rect 47068 19282 47124 19292
rect 47404 19010 47460 19022
rect 47404 18958 47406 19010
rect 47458 18958 47460 19010
rect 46620 18564 46676 18574
rect 46508 18562 46676 18564
rect 46508 18510 46622 18562
rect 46674 18510 46676 18562
rect 46508 18508 46676 18510
rect 46620 18498 46676 18508
rect 46956 18452 47012 18462
rect 46844 18450 47012 18452
rect 46844 18398 46958 18450
rect 47010 18398 47012 18450
rect 46844 18396 47012 18398
rect 46284 18274 46340 18284
rect 46732 18338 46788 18350
rect 46732 18286 46734 18338
rect 46786 18286 46788 18338
rect 46620 17780 46676 17790
rect 46732 17780 46788 18286
rect 46620 17778 46788 17780
rect 46620 17726 46622 17778
rect 46674 17726 46788 17778
rect 46620 17724 46788 17726
rect 46620 17714 46676 17724
rect 46844 17108 46900 18396
rect 46956 18386 47012 18396
rect 47404 17220 47460 18958
rect 47404 17154 47460 17164
rect 46172 15474 46228 15484
rect 46508 17052 46900 17108
rect 46508 15538 46564 17052
rect 46844 16884 46900 16894
rect 46508 15486 46510 15538
rect 46562 15486 46564 15538
rect 46284 15316 46340 15354
rect 46284 15250 46340 15260
rect 46508 15316 46564 15486
rect 46508 15250 46564 15260
rect 46620 16548 46676 16558
rect 46620 15148 46676 16492
rect 46620 15092 46788 15148
rect 46284 14532 46340 14542
rect 46732 14532 46788 15092
rect 46340 14476 46452 14532
rect 46284 14438 46340 14476
rect 46396 13970 46452 14476
rect 46396 13918 46398 13970
rect 46450 13918 46452 13970
rect 46396 13906 46452 13918
rect 46508 14476 46788 14532
rect 46508 14306 46564 14476
rect 46508 14254 46510 14306
rect 46562 14254 46564 14306
rect 46060 12350 46062 12402
rect 46114 12350 46116 12402
rect 45724 12180 45780 12190
rect 45388 11172 45444 11182
rect 45612 11172 45668 11182
rect 45388 11170 45556 11172
rect 45388 11118 45390 11170
rect 45442 11118 45556 11170
rect 45388 11116 45556 11118
rect 45388 11106 45444 11116
rect 45388 10612 45444 10622
rect 45388 10518 45444 10556
rect 44940 9998 44942 10050
rect 44994 9998 44996 10050
rect 44940 9986 44996 9998
rect 45052 9996 45332 10052
rect 45500 10052 45556 11116
rect 45612 11078 45668 11116
rect 45612 10836 45668 10846
rect 45724 10836 45780 12124
rect 46060 11788 46116 12350
rect 45836 11732 46116 11788
rect 46396 13748 46452 13758
rect 45836 11394 45892 11732
rect 45836 11342 45838 11394
rect 45890 11342 45892 11394
rect 45836 11330 45892 11342
rect 46284 11394 46340 11406
rect 46284 11342 46286 11394
rect 46338 11342 46340 11394
rect 45948 11284 46004 11294
rect 45948 11190 46004 11228
rect 46284 11172 46340 11342
rect 46284 11106 46340 11116
rect 45612 10834 45780 10836
rect 45612 10782 45614 10834
rect 45666 10782 45780 10834
rect 45612 10780 45780 10782
rect 45612 10770 45668 10780
rect 46396 10276 46452 13692
rect 46508 10836 46564 14254
rect 46844 14306 46900 16828
rect 47628 15092 47684 20972
rect 47740 20468 47796 21420
rect 47740 20412 48020 20468
rect 47852 19796 47908 19806
rect 47852 19702 47908 19740
rect 47964 19236 48020 20412
rect 48076 20020 48132 20030
rect 48076 19926 48132 19964
rect 48188 19236 48244 19246
rect 47964 19234 48244 19236
rect 47964 19182 48190 19234
rect 48242 19182 48244 19234
rect 47964 19180 48244 19182
rect 47740 19124 47796 19134
rect 47740 19030 47796 19068
rect 47852 18340 47908 18350
rect 48188 18340 48244 19180
rect 47852 18338 48244 18340
rect 47852 18286 47854 18338
rect 47906 18286 48244 18338
rect 47852 18284 48244 18286
rect 47852 17444 47908 18284
rect 47852 17378 47908 17388
rect 47628 15026 47684 15036
rect 48188 14530 48244 14542
rect 48188 14478 48190 14530
rect 48242 14478 48244 14530
rect 46844 14254 46846 14306
rect 46898 14254 46900 14306
rect 46844 13972 46900 14254
rect 46956 14418 47012 14430
rect 46956 14366 46958 14418
rect 47010 14366 47012 14418
rect 46956 14308 47012 14366
rect 47404 14308 47460 14318
rect 46956 14252 47404 14308
rect 47404 14214 47460 14252
rect 46844 13906 46900 13916
rect 46732 13858 46788 13870
rect 46732 13806 46734 13858
rect 46786 13806 46788 13858
rect 46732 13524 46788 13806
rect 46732 13458 46788 13468
rect 48188 13524 48244 14478
rect 48188 13458 48244 13468
rect 46956 11394 47012 11406
rect 46956 11342 46958 11394
rect 47010 11342 47012 11394
rect 46844 11284 46900 11294
rect 46956 11284 47012 11342
rect 46900 11228 47012 11284
rect 46844 11218 46900 11228
rect 46508 10780 46900 10836
rect 46396 10210 46452 10220
rect 46284 10164 46340 10174
rect 45500 9996 45780 10052
rect 44828 6692 44884 6702
rect 44828 6598 44884 6636
rect 44380 5170 44436 5180
rect 44492 5628 44772 5684
rect 44492 4564 44548 5628
rect 44940 5236 44996 5246
rect 44940 5142 44996 5180
rect 45052 5012 45108 9996
rect 45388 9828 45444 9838
rect 45164 9826 45444 9828
rect 45164 9774 45390 9826
rect 45442 9774 45444 9826
rect 45164 9772 45444 9774
rect 45164 9044 45220 9772
rect 45388 9762 45444 9772
rect 45612 9826 45668 9838
rect 45612 9774 45614 9826
rect 45666 9774 45668 9826
rect 45612 9380 45668 9774
rect 45388 9324 45668 9380
rect 45388 9044 45444 9324
rect 45164 9042 45332 9044
rect 45164 8990 45166 9042
rect 45218 8990 45332 9042
rect 45164 8988 45332 8990
rect 45164 8978 45220 8988
rect 45276 8428 45332 8988
rect 45388 8950 45444 8988
rect 45724 8930 45780 9996
rect 45836 9828 45892 9838
rect 45836 9826 46004 9828
rect 45836 9774 45838 9826
rect 45890 9774 46004 9826
rect 45836 9772 46004 9774
rect 45836 9762 45892 9772
rect 45948 9716 46004 9772
rect 45948 9650 46004 9660
rect 46060 9714 46116 9726
rect 46060 9662 46062 9714
rect 46114 9662 46116 9714
rect 45724 8878 45726 8930
rect 45778 8878 45780 8930
rect 45724 8866 45780 8878
rect 45836 9044 45892 9054
rect 46060 9044 46116 9662
rect 45836 9042 46116 9044
rect 45836 8990 45838 9042
rect 45890 8990 46116 9042
rect 45836 8988 46116 8990
rect 46172 9716 46228 9726
rect 45276 8372 45444 8428
rect 45388 7700 45444 8372
rect 45388 6802 45444 7644
rect 45388 6750 45390 6802
rect 45442 6750 45444 6802
rect 45388 6738 45444 6750
rect 45724 6692 45780 6702
rect 45836 6692 45892 8988
rect 45948 8820 46004 8830
rect 46172 8820 46228 9660
rect 46284 9604 46340 10108
rect 46396 9828 46452 9838
rect 46396 9734 46452 9772
rect 46844 9826 46900 10780
rect 47964 10612 48020 10622
rect 47404 10052 47460 10062
rect 47404 9958 47460 9996
rect 46844 9774 46846 9826
rect 46898 9774 46900 9826
rect 46844 9762 46900 9774
rect 47852 9828 47908 9838
rect 47852 9734 47908 9772
rect 46508 9604 46564 9614
rect 46284 9602 46564 9604
rect 46284 9550 46510 9602
rect 46562 9550 46564 9602
rect 46284 9548 46564 9550
rect 45948 8818 46228 8820
rect 45948 8766 45950 8818
rect 46002 8766 46228 8818
rect 45948 8764 46228 8766
rect 45948 8754 46004 8764
rect 45724 6690 46340 6692
rect 45724 6638 45726 6690
rect 45778 6638 46340 6690
rect 45724 6636 46340 6638
rect 45724 6580 45780 6636
rect 45724 6514 45780 6524
rect 46284 6578 46340 6636
rect 46284 6526 46286 6578
rect 46338 6526 46340 6578
rect 46284 6514 46340 6526
rect 46396 6468 46452 9548
rect 46508 9538 46564 9548
rect 47292 8484 47348 8494
rect 47292 8390 47348 8428
rect 46396 6402 46452 6412
rect 46508 8260 46564 8270
rect 46508 6690 46564 8204
rect 47180 8260 47236 8270
rect 47180 8166 47236 8204
rect 46732 7700 46788 7710
rect 47068 7700 47124 7710
rect 46788 7698 47124 7700
rect 46788 7646 47070 7698
rect 47122 7646 47124 7698
rect 46788 7644 47124 7646
rect 46732 7606 46788 7644
rect 47068 7634 47124 7644
rect 47740 7588 47796 7598
rect 46844 7476 46900 7486
rect 46844 7382 46900 7420
rect 47740 7474 47796 7532
rect 47740 7422 47742 7474
rect 47794 7422 47796 7474
rect 47740 7410 47796 7422
rect 47964 7476 48020 10556
rect 48076 9716 48132 9726
rect 48076 9622 48132 9660
rect 48188 9714 48244 9726
rect 48188 9662 48190 9714
rect 48242 9662 48244 9714
rect 48188 8260 48244 9662
rect 48300 9268 48356 23660
rect 48412 23380 48468 25230
rect 48412 23314 48468 23324
rect 48524 14308 48580 28028
rect 48636 27860 48692 33964
rect 48860 33926 48916 33964
rect 48748 33348 48804 33358
rect 48748 33254 48804 33292
rect 49084 33236 49140 34860
rect 49532 34850 49588 34860
rect 49756 34914 49812 35308
rect 49756 34862 49758 34914
rect 49810 34862 49812 34914
rect 49756 34850 49812 34862
rect 49868 35588 49924 35598
rect 49644 34804 49700 34814
rect 49644 34710 49700 34748
rect 49308 34692 49364 34702
rect 49196 34690 49364 34692
rect 49196 34638 49310 34690
rect 49362 34638 49364 34690
rect 49196 34636 49364 34638
rect 49196 34020 49252 34636
rect 49308 34626 49364 34636
rect 49756 34356 49812 34366
rect 49196 33954 49252 33964
rect 49644 34130 49700 34142
rect 49644 34078 49646 34130
rect 49698 34078 49700 34130
rect 49532 33796 49588 33806
rect 49420 33348 49476 33358
rect 49420 33254 49476 33292
rect 49084 33234 49364 33236
rect 49084 33182 49086 33234
rect 49138 33182 49364 33234
rect 49084 33180 49364 33182
rect 49084 33170 49140 33180
rect 49308 32786 49364 33180
rect 49308 32734 49310 32786
rect 49362 32734 49364 32786
rect 49308 32722 49364 32734
rect 49532 32788 49588 33740
rect 49644 33684 49700 34078
rect 49644 33618 49700 33628
rect 49756 33234 49812 34300
rect 49868 34244 49924 35532
rect 50092 34356 50148 36428
rect 50204 35308 50260 41132
rect 50876 41076 50932 42590
rect 50988 42866 51044 42878
rect 50988 42814 50990 42866
rect 51042 42814 51044 42866
rect 50988 42084 51044 42814
rect 51100 42084 51156 42094
rect 50988 42082 51156 42084
rect 50988 42030 51102 42082
rect 51154 42030 51156 42082
rect 50988 42028 51156 42030
rect 51100 42018 51156 42028
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50876 40628 50932 41020
rect 50764 40572 50932 40628
rect 50652 40402 50708 40414
rect 50652 40350 50654 40402
rect 50706 40350 50708 40402
rect 50428 39620 50484 39630
rect 50428 38836 50484 39564
rect 50540 39508 50596 39518
rect 50540 39414 50596 39452
rect 50652 39396 50708 40350
rect 50764 39506 50820 40572
rect 50876 39732 50932 39742
rect 50876 39730 51156 39732
rect 50876 39678 50878 39730
rect 50930 39678 51156 39730
rect 50876 39676 51156 39678
rect 50876 39666 50932 39676
rect 50764 39454 50766 39506
rect 50818 39454 50820 39506
rect 50764 39442 50820 39454
rect 50652 39330 50708 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 51100 38946 51156 39676
rect 51100 38894 51102 38946
rect 51154 38894 51156 38946
rect 51100 38882 51156 38894
rect 50428 38742 50484 38780
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50652 37266 50708 37278
rect 50652 37214 50654 37266
rect 50706 37214 50708 37266
rect 50652 36372 50708 37214
rect 50988 36484 51044 36494
rect 50988 36390 51044 36428
rect 51212 36484 51268 43484
rect 53004 43426 53060 43484
rect 53004 43374 53006 43426
rect 53058 43374 53060 43426
rect 53004 43362 53060 43374
rect 53228 42084 53284 42094
rect 53228 41858 53284 42028
rect 53228 41806 53230 41858
rect 53282 41806 53284 41858
rect 53228 41794 53284 41806
rect 51884 41298 51940 41310
rect 51884 41246 51886 41298
rect 51938 41246 51940 41298
rect 51884 40852 51940 41246
rect 51884 40786 51940 40796
rect 53004 40178 53060 40190
rect 53004 40126 53006 40178
rect 53058 40126 53060 40178
rect 53004 38164 53060 40126
rect 53228 39060 53284 39070
rect 53228 38722 53284 39004
rect 53228 38670 53230 38722
rect 53282 38670 53284 38722
rect 53228 38658 53284 38670
rect 53004 38098 53060 38108
rect 51212 36390 51268 36428
rect 53004 37042 53060 37054
rect 53004 36990 53006 37042
rect 53058 36990 53060 37042
rect 50652 36306 50708 36316
rect 50764 36260 50820 36298
rect 50764 36194 50820 36204
rect 51100 36258 51156 36270
rect 51100 36206 51102 36258
rect 51154 36206 51156 36258
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50316 35924 50372 35934
rect 50316 35698 50372 35868
rect 51100 35812 51156 36206
rect 50316 35646 50318 35698
rect 50370 35646 50372 35698
rect 50316 35634 50372 35646
rect 50876 35756 51156 35812
rect 50204 35252 50372 35308
rect 50092 34262 50148 34300
rect 49868 34178 49924 34188
rect 50316 34132 50372 35252
rect 50876 35138 50932 35756
rect 50876 35086 50878 35138
rect 50930 35086 50932 35138
rect 50876 35074 50932 35086
rect 51100 35586 51156 35598
rect 51100 35534 51102 35586
rect 51154 35534 51156 35586
rect 51100 35026 51156 35534
rect 53004 35476 53060 36990
rect 53228 36484 53284 36494
rect 53228 35586 53284 36428
rect 53228 35534 53230 35586
rect 53282 35534 53284 35586
rect 53228 35522 53284 35534
rect 53004 35410 53060 35420
rect 51100 34974 51102 35026
rect 51154 34974 51156 35026
rect 51100 34962 51156 34974
rect 50652 34692 50708 34702
rect 51100 34692 51156 34702
rect 50652 34690 51156 34692
rect 50652 34638 50654 34690
rect 50706 34638 51102 34690
rect 51154 34638 51156 34690
rect 50652 34636 51156 34638
rect 50652 34626 50708 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 34130 50484 34132
rect 50316 34078 50318 34130
rect 50370 34078 50484 34130
rect 50316 34076 50484 34078
rect 50316 34066 50372 34076
rect 50204 34020 50260 34030
rect 50204 33926 50260 33964
rect 49756 33182 49758 33234
rect 49810 33182 49812 33234
rect 49756 33170 49812 33182
rect 50092 33908 50148 33918
rect 50092 33012 50148 33852
rect 50204 33122 50260 33134
rect 50204 33070 50206 33122
rect 50258 33070 50260 33122
rect 50204 33012 50260 33070
rect 49980 32956 50260 33012
rect 49868 32788 49924 32798
rect 49532 32786 49924 32788
rect 49532 32734 49534 32786
rect 49586 32734 49870 32786
rect 49922 32734 49924 32786
rect 49532 32732 49924 32734
rect 49532 32722 49588 32732
rect 49868 32722 49924 32732
rect 49084 32452 49140 32462
rect 49084 32358 49140 32396
rect 49420 32450 49476 32462
rect 49420 32398 49422 32450
rect 49474 32398 49476 32450
rect 48860 32340 48916 32350
rect 49420 32340 49476 32398
rect 49756 32340 49812 32350
rect 49420 32338 49812 32340
rect 49420 32286 49758 32338
rect 49810 32286 49812 32338
rect 49420 32284 49812 32286
rect 48860 32246 48916 32284
rect 49756 32274 49812 32284
rect 48972 31554 49028 31566
rect 48972 31502 48974 31554
rect 49026 31502 49028 31554
rect 48972 30884 49028 31502
rect 49868 31556 49924 31566
rect 49868 31462 49924 31500
rect 48972 30818 49028 30828
rect 49980 30884 50036 32956
rect 50092 32788 50148 32798
rect 50092 32786 50260 32788
rect 50092 32734 50094 32786
rect 50146 32734 50260 32786
rect 50092 32732 50260 32734
rect 50092 32722 50148 32732
rect 50092 32338 50148 32350
rect 50092 32286 50094 32338
rect 50146 32286 50148 32338
rect 50092 32004 50148 32286
rect 50204 32228 50260 32732
rect 50316 32452 50372 32462
rect 50428 32452 50484 34076
rect 50652 34130 50708 34142
rect 50652 34078 50654 34130
rect 50706 34078 50708 34130
rect 50652 33796 50708 34078
rect 50652 33730 50708 33740
rect 50876 34020 50932 34030
rect 50876 33570 50932 33964
rect 50876 33518 50878 33570
rect 50930 33518 50932 33570
rect 50876 33506 50932 33518
rect 50988 33124 51044 33134
rect 50988 33030 51044 33068
rect 51100 33124 51156 34636
rect 53004 33906 53060 33918
rect 53004 33854 53006 33906
rect 53058 33854 53060 33906
rect 51660 33124 51716 33134
rect 51100 33122 51716 33124
rect 51100 33070 51102 33122
rect 51154 33070 51662 33122
rect 51714 33070 51716 33122
rect 51100 33068 51716 33070
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50316 32450 50484 32452
rect 50316 32398 50318 32450
rect 50370 32398 50484 32450
rect 50316 32396 50484 32398
rect 50316 32386 50372 32396
rect 50204 32172 50372 32228
rect 50204 32004 50260 32014
rect 50092 32002 50260 32004
rect 50092 31950 50206 32002
rect 50258 31950 50260 32002
rect 50092 31948 50260 31950
rect 50204 31938 50260 31948
rect 49644 30324 49700 30334
rect 49084 29314 49140 29326
rect 49084 29262 49086 29314
rect 49138 29262 49140 29314
rect 49084 28868 49140 29262
rect 49084 28802 49140 28812
rect 48972 28756 49028 28766
rect 48636 27794 48692 27804
rect 48748 28418 48804 28430
rect 48748 28366 48750 28418
rect 48802 28366 48804 28418
rect 48748 26908 48804 28366
rect 48972 28082 49028 28700
rect 49084 28644 49140 28654
rect 49084 28550 49140 28588
rect 49644 28642 49700 30268
rect 49644 28590 49646 28642
rect 49698 28590 49700 28642
rect 48972 28030 48974 28082
rect 49026 28030 49028 28082
rect 48972 28018 49028 28030
rect 49644 26908 49700 28590
rect 49980 29428 50036 30828
rect 50316 30882 50372 32172
rect 50540 31892 50596 31902
rect 50540 31798 50596 31836
rect 50316 30830 50318 30882
rect 50370 30830 50372 30882
rect 50316 30818 50372 30830
rect 50428 31556 50484 31566
rect 50428 30324 50484 31500
rect 51100 31556 51156 33068
rect 51660 33058 51716 33068
rect 52444 33124 52500 33134
rect 52444 32674 52500 33068
rect 53004 32788 53060 33854
rect 53004 32722 53060 32732
rect 52444 32622 52446 32674
rect 52498 32622 52500 32674
rect 52444 32610 52500 32622
rect 53116 32562 53172 32574
rect 53116 32510 53118 32562
rect 53170 32510 53172 32562
rect 51100 31490 51156 31500
rect 52444 31892 52500 31902
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 52444 31106 52500 31836
rect 52444 31054 52446 31106
rect 52498 31054 52500 31106
rect 52444 31042 52500 31054
rect 53116 30994 53172 32510
rect 53116 30942 53118 30994
rect 53170 30942 53172 30994
rect 49980 27748 50036 29372
rect 49980 27654 50036 27692
rect 50092 30268 50484 30324
rect 52892 30324 52948 30334
rect 48748 26852 49028 26908
rect 48860 24834 48916 24846
rect 48860 24782 48862 24834
rect 48914 24782 48916 24834
rect 48748 24724 48804 24734
rect 48748 23380 48804 24668
rect 48860 24612 48916 24782
rect 48860 24546 48916 24556
rect 48748 23324 48916 23380
rect 48748 23156 48804 23166
rect 48748 23062 48804 23100
rect 48860 22932 48916 23324
rect 48748 22876 48916 22932
rect 48748 20020 48804 22876
rect 48636 19964 48804 20020
rect 48860 20130 48916 20142
rect 48860 20078 48862 20130
rect 48914 20078 48916 20130
rect 48636 19572 48692 19964
rect 48748 19796 48804 19806
rect 48748 19702 48804 19740
rect 48636 19516 48804 19572
rect 48636 18340 48692 18350
rect 48636 16098 48692 18284
rect 48748 18228 48804 19516
rect 48748 18162 48804 18172
rect 48748 17780 48804 17790
rect 48860 17780 48916 20078
rect 48748 17778 48916 17780
rect 48748 17726 48750 17778
rect 48802 17726 48916 17778
rect 48748 17724 48916 17726
rect 48748 17714 48804 17724
rect 48636 16046 48638 16098
rect 48690 16046 48692 16098
rect 48636 15204 48692 16046
rect 48860 16098 48916 17724
rect 48860 16046 48862 16098
rect 48914 16046 48916 16098
rect 48860 16034 48916 16046
rect 48748 15874 48804 15886
rect 48748 15822 48750 15874
rect 48802 15822 48804 15874
rect 48748 15426 48804 15822
rect 48972 15652 49028 26852
rect 49196 26852 49700 26908
rect 49196 26514 49252 26852
rect 49196 26462 49198 26514
rect 49250 26462 49252 26514
rect 49196 26450 49252 26462
rect 49868 26404 49924 26414
rect 49868 26310 49924 26348
rect 49084 26292 49140 26302
rect 49756 26292 49812 26302
rect 49084 26290 49812 26292
rect 49084 26238 49086 26290
rect 49138 26238 49758 26290
rect 49810 26238 49812 26290
rect 49084 26236 49812 26238
rect 49084 26226 49140 26236
rect 49196 26066 49252 26078
rect 49196 26014 49198 26066
rect 49250 26014 49252 26066
rect 49196 25506 49252 26014
rect 49196 25454 49198 25506
rect 49250 25454 49252 25506
rect 49196 25442 49252 25454
rect 49532 25396 49588 25406
rect 49532 25282 49588 25340
rect 49532 25230 49534 25282
rect 49586 25230 49588 25282
rect 49532 25218 49588 25230
rect 49644 25394 49700 25406
rect 49644 25342 49646 25394
rect 49698 25342 49700 25394
rect 49644 25060 49700 25342
rect 49084 25004 49700 25060
rect 49084 24946 49140 25004
rect 49756 24948 49812 26236
rect 49868 26068 49924 26078
rect 49868 25974 49924 26012
rect 49868 25508 49924 25518
rect 49868 25414 49924 25452
rect 49084 24894 49086 24946
rect 49138 24894 49140 24946
rect 49084 24882 49140 24894
rect 49644 24892 49812 24948
rect 49420 24724 49476 24734
rect 49420 24630 49476 24668
rect 49308 23716 49364 23726
rect 49196 23380 49252 23390
rect 49196 22484 49252 23324
rect 49308 23378 49364 23660
rect 49308 23326 49310 23378
rect 49362 23326 49364 23378
rect 49308 23314 49364 23326
rect 49644 23154 49700 24892
rect 49868 24724 49924 24734
rect 49868 24050 49924 24668
rect 49868 23998 49870 24050
rect 49922 23998 49924 24050
rect 49868 23940 49924 23998
rect 50092 23940 50148 30268
rect 52892 30098 52948 30268
rect 52892 30046 52894 30098
rect 52946 30046 52948 30098
rect 52892 30034 52948 30046
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 51212 29540 51268 29550
rect 51212 29446 51268 29484
rect 51884 29428 51940 29438
rect 51884 29334 51940 29372
rect 52444 29428 52500 29438
rect 52444 29334 52500 29372
rect 53116 29428 53172 30942
rect 53228 30100 53284 30110
rect 53284 30044 53396 30100
rect 53228 30006 53284 30044
rect 53340 29650 53396 30044
rect 53340 29598 53342 29650
rect 53394 29598 53396 29650
rect 53340 29586 53396 29598
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 53116 27858 53172 29372
rect 53116 27806 53118 27858
rect 53170 27806 53172 27858
rect 53116 27794 53172 27806
rect 50316 27746 50372 27758
rect 50316 27694 50318 27746
rect 50370 27694 50372 27746
rect 50316 25508 50372 27694
rect 52444 27746 52500 27758
rect 52444 27694 52446 27746
rect 52498 27694 52500 27746
rect 51660 27300 51716 27310
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 51660 26514 51716 27244
rect 52444 27300 52500 27694
rect 52444 27234 52500 27244
rect 53340 27412 53396 27422
rect 53228 27076 53284 27086
rect 53340 27076 53396 27356
rect 53228 27074 53396 27076
rect 53228 27022 53230 27074
rect 53282 27022 53396 27074
rect 53228 27020 53396 27022
rect 53228 27010 53284 27020
rect 51660 26462 51662 26514
rect 51714 26462 51716 26514
rect 51660 26450 51716 26462
rect 52892 26962 52948 26974
rect 52892 26910 52894 26962
rect 52946 26910 52948 26962
rect 52892 26404 52948 26910
rect 53340 26514 53396 27020
rect 53340 26462 53342 26514
rect 53394 26462 53396 26514
rect 53340 26450 53396 26462
rect 52892 26338 52948 26348
rect 51212 26292 51268 26302
rect 51884 26292 51940 26302
rect 51212 26290 52052 26292
rect 51212 26238 51214 26290
rect 51266 26238 51886 26290
rect 51938 26238 52052 26290
rect 51212 26236 52052 26238
rect 51212 26226 51268 26236
rect 51884 26226 51940 26236
rect 51548 26068 51604 26078
rect 51436 26066 51604 26068
rect 51436 26014 51550 26066
rect 51602 26014 51604 26066
rect 51436 26012 51604 26014
rect 50316 25452 50484 25508
rect 50204 25396 50260 25406
rect 50204 25302 50260 25340
rect 50428 25394 50484 25452
rect 50428 25342 50430 25394
rect 50482 25342 50484 25394
rect 50428 24948 50484 25342
rect 50876 25506 50932 25518
rect 50876 25454 50878 25506
rect 50930 25454 50932 25506
rect 50540 25284 50596 25322
rect 50540 25218 50596 25228
rect 50876 25172 50932 25454
rect 51100 25508 51156 25518
rect 51100 25414 51156 25452
rect 51324 25394 51380 25406
rect 51324 25342 51326 25394
rect 51378 25342 51380 25394
rect 51324 25172 51380 25342
rect 50556 25116 50820 25126
rect 50876 25116 51268 25172
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50652 24948 50708 24958
rect 50428 24946 50708 24948
rect 50428 24894 50654 24946
rect 50706 24894 50708 24946
rect 50428 24892 50708 24894
rect 50652 24882 50708 24892
rect 50764 24948 50820 24958
rect 50316 24724 50372 24734
rect 50204 24612 50260 24622
rect 50204 24518 50260 24556
rect 50092 23884 50260 23940
rect 49868 23874 49924 23884
rect 49756 23716 49812 23726
rect 49756 23378 49812 23660
rect 49756 23326 49758 23378
rect 49810 23326 49812 23378
rect 49756 23314 49812 23326
rect 50092 23714 50148 23726
rect 50092 23662 50094 23714
rect 50146 23662 50148 23714
rect 49644 23102 49646 23154
rect 49698 23102 49700 23154
rect 49644 22932 49700 23102
rect 49196 22390 49252 22428
rect 49308 22876 49700 22932
rect 49756 22930 49812 22942
rect 49756 22878 49758 22930
rect 49810 22878 49812 22930
rect 49084 19796 49140 19806
rect 49308 19796 49364 22876
rect 49756 21586 49812 22878
rect 49980 22260 50036 22270
rect 49980 21810 50036 22204
rect 49980 21758 49982 21810
rect 50034 21758 50036 21810
rect 49980 21746 50036 21758
rect 49756 21534 49758 21586
rect 49810 21534 49812 21586
rect 49756 21522 49812 21534
rect 50092 21586 50148 23662
rect 50092 21534 50094 21586
rect 50146 21534 50148 21586
rect 50092 21522 50148 21534
rect 49532 20580 49588 20590
rect 49084 19794 49364 19796
rect 49084 19742 49086 19794
rect 49138 19742 49364 19794
rect 49084 19740 49364 19742
rect 49420 20578 49588 20580
rect 49420 20526 49534 20578
rect 49586 20526 49588 20578
rect 49420 20524 49588 20526
rect 49420 20018 49476 20524
rect 49532 20514 49588 20524
rect 49868 20580 49924 20590
rect 49868 20486 49924 20524
rect 49420 19966 49422 20018
rect 49474 19966 49476 20018
rect 49084 19124 49140 19740
rect 49308 19348 49364 19358
rect 49084 19058 49140 19068
rect 49196 19292 49308 19348
rect 49196 17668 49252 19292
rect 49308 19254 49364 19292
rect 49084 17612 49196 17668
rect 49084 15764 49140 17612
rect 49196 17574 49252 17612
rect 49420 18450 49476 19966
rect 49756 20130 49812 20142
rect 49756 20078 49758 20130
rect 49810 20078 49812 20130
rect 49756 20020 49812 20078
rect 49756 19954 49812 19964
rect 49420 18398 49422 18450
rect 49474 18398 49476 18450
rect 49196 17444 49252 17454
rect 49196 16882 49252 17388
rect 49308 16996 49364 17006
rect 49308 16902 49364 16940
rect 49196 16830 49198 16882
rect 49250 16830 49252 16882
rect 49196 16548 49252 16830
rect 49420 16772 49476 18398
rect 49644 18562 49700 18574
rect 49644 18510 49646 18562
rect 49698 18510 49700 18562
rect 49644 18340 49700 18510
rect 49644 18274 49700 18284
rect 49196 16482 49252 16492
rect 49308 16716 49476 16772
rect 49532 16882 49588 16894
rect 49532 16830 49534 16882
rect 49586 16830 49588 16882
rect 49196 15988 49252 15998
rect 49196 15894 49252 15932
rect 49084 15708 49252 15764
rect 48972 15596 49140 15652
rect 49084 15540 49140 15596
rect 49084 15474 49140 15484
rect 48748 15374 48750 15426
rect 48802 15374 48804 15426
rect 48748 15362 48804 15374
rect 49084 15316 49140 15326
rect 49084 15222 49140 15260
rect 48636 15138 48692 15148
rect 48860 15202 48916 15214
rect 48860 15150 48862 15202
rect 48914 15150 48916 15202
rect 48860 14642 48916 15150
rect 48860 14590 48862 14642
rect 48914 14590 48916 14642
rect 48860 14578 48916 14590
rect 48524 14242 48580 14252
rect 49196 13524 49252 15708
rect 49196 13458 49252 13468
rect 49308 12628 49364 16716
rect 49532 16098 49588 16830
rect 49532 16046 49534 16098
rect 49586 16046 49588 16098
rect 49532 16034 49588 16046
rect 50092 16098 50148 16110
rect 50092 16046 50094 16098
rect 50146 16046 50148 16098
rect 49756 15988 49812 15998
rect 49756 15894 49812 15932
rect 49980 15988 50036 15998
rect 49980 15894 50036 15932
rect 49084 12572 49364 12628
rect 49644 15540 49700 15550
rect 49084 12180 49140 12572
rect 49644 12516 49700 15484
rect 50092 15428 50148 16046
rect 50092 15148 50148 15372
rect 49084 12114 49140 12124
rect 49308 12460 49700 12516
rect 49868 15092 50148 15148
rect 49196 12066 49252 12078
rect 49196 12014 49198 12066
rect 49250 12014 49252 12066
rect 49084 11506 49140 11518
rect 49084 11454 49086 11506
rect 49138 11454 49140 11506
rect 48300 9202 48356 9212
rect 48412 9826 48468 9838
rect 48412 9774 48414 9826
rect 48466 9774 48468 9826
rect 48188 8194 48244 8204
rect 48300 7588 48356 7598
rect 47964 7474 48244 7476
rect 47964 7422 47966 7474
rect 48018 7422 48244 7474
rect 47964 7420 48244 7422
rect 47964 7410 48020 7420
rect 46508 6638 46510 6690
rect 46562 6638 46564 6690
rect 45164 5012 45220 5022
rect 45052 4956 45164 5012
rect 45164 4946 45220 4956
rect 44828 4900 44884 4910
rect 44492 4470 44548 4508
rect 44604 4898 44884 4900
rect 44604 4846 44830 4898
rect 44882 4846 44884 4898
rect 44604 4844 44884 4846
rect 44604 4116 44660 4844
rect 44828 4834 44884 4844
rect 44380 4060 44660 4116
rect 44380 3666 44436 4060
rect 44380 3614 44382 3666
rect 44434 3614 44436 3666
rect 44380 3602 44436 3614
rect 46508 3666 46564 6638
rect 46732 7250 46788 7262
rect 46732 7198 46734 7250
rect 46786 7198 46788 7250
rect 46732 6692 46788 7198
rect 47516 7250 47572 7262
rect 47516 7198 47518 7250
rect 47570 7198 47572 7250
rect 47516 6916 47572 7198
rect 47516 6860 48020 6916
rect 46732 6626 46788 6636
rect 47404 6692 47460 6702
rect 47404 6598 47460 6636
rect 47628 6692 47684 6702
rect 47628 6598 47684 6636
rect 47852 6690 47908 6702
rect 47852 6638 47854 6690
rect 47906 6638 47908 6690
rect 47180 6580 47236 6590
rect 47180 6486 47236 6524
rect 47628 6466 47684 6478
rect 47628 6414 47630 6466
rect 47682 6414 47684 6466
rect 46732 5124 46788 5134
rect 46732 5030 46788 5068
rect 47404 5010 47460 5022
rect 47404 4958 47406 5010
rect 47458 4958 47460 5010
rect 47404 4564 47460 4958
rect 47516 4564 47572 4574
rect 47404 4562 47572 4564
rect 47404 4510 47518 4562
rect 47570 4510 47572 4562
rect 47404 4508 47572 4510
rect 47516 4498 47572 4508
rect 47628 4450 47684 6414
rect 47852 6468 47908 6638
rect 47964 6692 48020 6860
rect 48076 6692 48132 6702
rect 47964 6636 48076 6692
rect 48076 6598 48132 6636
rect 48188 6580 48244 7420
rect 48300 6692 48356 7532
rect 48412 7028 48468 9774
rect 49084 9716 49140 11454
rect 49196 11172 49252 12014
rect 49196 11106 49252 11116
rect 49196 10610 49252 10622
rect 49196 10558 49198 10610
rect 49250 10558 49252 10610
rect 49196 10164 49252 10558
rect 49196 10098 49252 10108
rect 49084 8258 49140 9660
rect 49084 8206 49086 8258
rect 49138 8206 49140 8258
rect 49084 8194 49140 8206
rect 48636 8146 48692 8158
rect 48636 8094 48638 8146
rect 48690 8094 48692 8146
rect 48412 6962 48468 6972
rect 48524 7476 48580 7486
rect 48524 6802 48580 7420
rect 48524 6750 48526 6802
rect 48578 6750 48580 6802
rect 48524 6738 48580 6750
rect 48412 6692 48468 6702
rect 48300 6690 48468 6692
rect 48300 6638 48414 6690
rect 48466 6638 48468 6690
rect 48300 6636 48468 6638
rect 48412 6626 48468 6636
rect 48636 6692 48692 8094
rect 49308 7140 49364 12460
rect 49868 12404 49924 15092
rect 50204 14644 50260 23884
rect 50316 23826 50372 24668
rect 50540 24722 50596 24734
rect 50764 24724 50820 24892
rect 50876 24836 50932 24846
rect 50876 24742 50932 24780
rect 50540 24670 50542 24722
rect 50594 24670 50596 24722
rect 50428 23940 50484 23950
rect 50540 23940 50596 24670
rect 50484 23884 50596 23940
rect 50652 24668 50820 24724
rect 51212 24724 51268 25116
rect 51324 25106 51380 25116
rect 51436 24948 51492 26012
rect 51548 26002 51604 26012
rect 51660 26068 51716 26078
rect 51660 25506 51716 26012
rect 51660 25454 51662 25506
rect 51714 25454 51716 25506
rect 51660 25442 51716 25454
rect 51548 25282 51604 25294
rect 51548 25230 51550 25282
rect 51602 25230 51604 25282
rect 51548 25172 51604 25230
rect 51548 25116 51940 25172
rect 51548 24948 51604 24958
rect 51436 24946 51604 24948
rect 51436 24894 51550 24946
rect 51602 24894 51604 24946
rect 51436 24892 51604 24894
rect 51548 24882 51604 24892
rect 51436 24724 51492 24734
rect 51660 24724 51716 24734
rect 51212 24722 51604 24724
rect 51212 24670 51438 24722
rect 51490 24670 51604 24722
rect 51212 24668 51604 24670
rect 50428 23846 50484 23884
rect 50316 23774 50318 23826
rect 50370 23774 50372 23826
rect 50316 23042 50372 23774
rect 50652 23716 50708 24668
rect 51436 24658 51492 24668
rect 50316 22990 50318 23042
rect 50370 22990 50372 23042
rect 50316 22978 50372 22990
rect 50428 23660 50708 23716
rect 50876 23714 50932 23726
rect 50876 23662 50878 23714
rect 50930 23662 50932 23714
rect 50428 21698 50484 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50876 23156 50932 23662
rect 50876 23090 50932 23100
rect 51324 22370 51380 22382
rect 51324 22318 51326 22370
rect 51378 22318 51380 22370
rect 50988 22260 51044 22270
rect 50988 22166 51044 22204
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50428 21646 50430 21698
rect 50482 21646 50484 21698
rect 50428 20804 50484 21646
rect 50316 20748 50484 20804
rect 50316 20244 50372 20748
rect 50316 20178 50372 20188
rect 50428 20578 50484 20590
rect 50428 20526 50430 20578
rect 50482 20526 50484 20578
rect 50316 20020 50372 20030
rect 50428 20020 50484 20526
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 20018 50484 20020
rect 50316 19966 50318 20018
rect 50370 19966 50484 20018
rect 50316 19964 50484 19966
rect 50316 19348 50372 19964
rect 50316 19282 50372 19292
rect 51100 19906 51156 19918
rect 51100 19854 51102 19906
rect 51154 19854 51156 19906
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50988 18676 51044 18686
rect 51100 18676 51156 19854
rect 51324 19908 51380 22318
rect 51436 22260 51492 22270
rect 51436 22166 51492 22204
rect 51548 22258 51604 24668
rect 51660 24630 51716 24668
rect 51884 24722 51940 25116
rect 51884 24670 51886 24722
rect 51938 24670 51940 24722
rect 51884 24658 51940 24670
rect 51996 23828 52052 26236
rect 53228 25394 53284 25406
rect 53228 25342 53230 25394
rect 53282 25342 53284 25394
rect 52892 25282 52948 25294
rect 52892 25230 52894 25282
rect 52946 25230 52948 25282
rect 52108 23828 52164 23838
rect 51996 23772 52108 23828
rect 51548 22206 51550 22258
rect 51602 22206 51604 22258
rect 51324 19842 51380 19852
rect 51548 20580 51604 22206
rect 52108 22146 52164 23772
rect 52892 23716 52948 25230
rect 53228 24724 53284 25342
rect 53228 24630 53284 24668
rect 52892 23650 52948 23660
rect 53116 23156 53172 23166
rect 53116 23062 53172 23100
rect 52444 23044 52500 23054
rect 52444 23042 52836 23044
rect 52444 22990 52446 23042
rect 52498 22990 52836 23042
rect 52444 22988 52836 22990
rect 52444 22978 52500 22988
rect 52780 22482 52836 22988
rect 52780 22430 52782 22482
rect 52834 22430 52836 22482
rect 52780 22418 52836 22430
rect 52668 22260 52724 22270
rect 52668 22166 52724 22204
rect 52108 22094 52110 22146
rect 52162 22094 52164 22146
rect 52108 22036 52164 22094
rect 52892 22146 52948 22158
rect 52892 22094 52894 22146
rect 52946 22094 52948 22146
rect 52892 22036 52948 22094
rect 52108 21980 52948 22036
rect 53228 22036 53284 22046
rect 52668 21700 52724 21710
rect 52668 21606 52724 21644
rect 52892 21700 52948 21710
rect 53228 21700 53284 21980
rect 52892 21698 53060 21700
rect 52892 21646 52894 21698
rect 52946 21646 53060 21698
rect 52892 21644 53060 21646
rect 52892 21634 52948 21644
rect 50988 18674 51156 18676
rect 50988 18622 50990 18674
rect 51042 18622 51156 18674
rect 50988 18620 51156 18622
rect 50988 18610 51044 18620
rect 51436 18564 51492 18574
rect 51548 18564 51604 20524
rect 51772 19908 51828 19918
rect 51436 18562 51604 18564
rect 51436 18510 51438 18562
rect 51490 18510 51604 18562
rect 51436 18508 51604 18510
rect 51660 19852 51772 19908
rect 51436 18498 51492 18508
rect 50764 18452 50820 18462
rect 50428 18450 50820 18452
rect 50428 18398 50766 18450
rect 50818 18398 50820 18450
rect 50428 18396 50820 18398
rect 50428 16772 50484 18396
rect 50764 18386 50820 18396
rect 50988 18452 51044 18462
rect 50988 17668 51044 18396
rect 51548 18338 51604 18350
rect 51548 18286 51550 18338
rect 51602 18286 51604 18338
rect 51100 18228 51156 18238
rect 51548 18228 51604 18286
rect 51100 18226 51604 18228
rect 51100 18174 51102 18226
rect 51154 18174 51604 18226
rect 51100 18172 51604 18174
rect 51100 18162 51156 18172
rect 51212 18004 51268 18014
rect 51212 17890 51268 17948
rect 51212 17838 51214 17890
rect 51266 17838 51268 17890
rect 51212 17826 51268 17838
rect 51660 17780 51716 19852
rect 51772 19842 51828 19852
rect 52220 19348 52276 19358
rect 52220 19254 52276 19292
rect 52892 19012 52948 19022
rect 52780 19010 52948 19012
rect 52780 18958 52894 19010
rect 52946 18958 52948 19010
rect 52780 18956 52948 18958
rect 51772 18450 51828 18462
rect 51772 18398 51774 18450
rect 51826 18398 51828 18450
rect 51772 18004 51828 18398
rect 51884 18452 51940 18462
rect 51884 18358 51940 18396
rect 52220 18450 52276 18462
rect 52220 18398 52222 18450
rect 52274 18398 52276 18450
rect 52220 18228 52276 18398
rect 52444 18452 52500 18462
rect 52444 18358 52500 18396
rect 52556 18450 52612 18462
rect 52556 18398 52558 18450
rect 52610 18398 52612 18450
rect 52220 18162 52276 18172
rect 51772 17938 51828 17948
rect 52108 18004 52164 18014
rect 51660 17724 51828 17780
rect 50988 17602 51044 17612
rect 51212 17668 51268 17678
rect 50540 17554 50596 17566
rect 50540 17502 50542 17554
rect 50594 17502 50596 17554
rect 50540 17444 50596 17502
rect 50652 17556 50708 17566
rect 50652 17462 50708 17500
rect 51100 17554 51156 17566
rect 51100 17502 51102 17554
rect 51154 17502 51156 17554
rect 50540 17378 50596 17388
rect 50876 17442 50932 17454
rect 50876 17390 50878 17442
rect 50930 17390 50932 17442
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50316 16716 50484 16772
rect 50316 15540 50372 16716
rect 50876 16436 50932 17390
rect 51100 17444 51156 17502
rect 51212 17554 51268 17612
rect 51212 17502 51214 17554
rect 51266 17502 51268 17554
rect 51212 17490 51268 17502
rect 51660 17554 51716 17566
rect 51660 17502 51662 17554
rect 51714 17502 51716 17554
rect 51100 17378 51156 17388
rect 50876 16370 50932 16380
rect 51324 17108 51380 17118
rect 51660 17108 51716 17502
rect 51772 17554 51828 17724
rect 51996 17666 52052 17678
rect 51996 17614 51998 17666
rect 52050 17614 52052 17666
rect 51996 17556 52052 17614
rect 51772 17502 51774 17554
rect 51826 17502 51828 17554
rect 51772 17490 51828 17502
rect 51884 17500 52052 17556
rect 51884 17444 51940 17500
rect 51884 17378 51940 17388
rect 51772 17108 51828 17118
rect 51660 17052 51772 17108
rect 51828 17052 51940 17108
rect 51212 16212 51268 16222
rect 51324 16212 51380 17052
rect 51772 17014 51828 17052
rect 50764 16210 51380 16212
rect 50764 16158 51214 16210
rect 51266 16158 51380 16210
rect 50764 16156 51380 16158
rect 51548 16660 51604 16670
rect 50764 16098 50820 16156
rect 51212 16146 51268 16156
rect 50764 16046 50766 16098
rect 50818 16046 50820 16098
rect 50764 16034 50820 16046
rect 50428 15988 50484 15998
rect 50428 15894 50484 15932
rect 50652 15876 50708 15914
rect 50652 15810 50708 15820
rect 51324 15876 51380 15886
rect 51380 15820 51492 15876
rect 51324 15810 51380 15820
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50316 15474 50372 15484
rect 51100 15316 51156 15326
rect 51100 15222 51156 15260
rect 51436 15314 51492 15820
rect 51436 15262 51438 15314
rect 51490 15262 51492 15314
rect 51324 15204 51380 15242
rect 51324 15138 51380 15148
rect 51436 14868 51492 15262
rect 50204 14578 50260 14588
rect 50988 14812 51492 14868
rect 50988 14642 51044 14812
rect 50988 14590 50990 14642
rect 51042 14590 51044 14642
rect 50988 14578 51044 14590
rect 51436 14306 51492 14318
rect 51436 14254 51438 14306
rect 51490 14254 51492 14306
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51100 13524 51156 13534
rect 49420 12402 49924 12404
rect 49420 12350 49870 12402
rect 49922 12350 49924 12402
rect 49420 12348 49924 12350
rect 49420 10836 49476 12348
rect 49868 12338 49924 12348
rect 50316 13412 50372 13422
rect 49532 12180 49588 12190
rect 49532 12086 49588 12124
rect 50316 12178 50372 13356
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 51100 12290 51156 13468
rect 51436 13412 51492 14254
rect 51436 13346 51492 13356
rect 51100 12238 51102 12290
rect 51154 12238 51156 12290
rect 51100 12226 51156 12238
rect 50316 12126 50318 12178
rect 50370 12126 50372 12178
rect 49532 11172 49588 11182
rect 49980 11172 50036 11182
rect 49588 11170 50036 11172
rect 49588 11118 49982 11170
rect 50034 11118 50036 11170
rect 49588 11116 50036 11118
rect 49532 11078 49588 11116
rect 49644 10836 49700 10846
rect 49420 10780 49588 10836
rect 49420 10612 49476 10622
rect 49532 10612 49588 10780
rect 49644 10742 49700 10780
rect 49644 10612 49700 10622
rect 49532 10610 49700 10612
rect 49532 10558 49646 10610
rect 49698 10558 49700 10610
rect 49532 10556 49700 10558
rect 49420 9716 49476 10556
rect 49644 10546 49700 10556
rect 49868 10610 49924 10622
rect 49868 10558 49870 10610
rect 49922 10558 49924 10610
rect 49868 9940 49924 10558
rect 49980 10612 50036 11116
rect 50316 10612 50372 12126
rect 50652 11282 50708 11294
rect 50652 11230 50654 11282
rect 50706 11230 50708 11282
rect 50652 11172 50708 11230
rect 50652 11106 50708 11116
rect 50764 11172 50820 11182
rect 50764 11170 51156 11172
rect 50764 11118 50766 11170
rect 50818 11118 51156 11170
rect 50764 11116 51156 11118
rect 50764 11106 50820 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 51100 10722 51156 11116
rect 51100 10670 51102 10722
rect 51154 10670 51156 10722
rect 51100 10658 51156 10670
rect 49980 10610 50372 10612
rect 49980 10558 50318 10610
rect 50370 10558 50372 10610
rect 49980 10556 50372 10558
rect 49868 9884 50036 9940
rect 49756 9828 49812 9838
rect 49532 9716 49588 9726
rect 49420 9714 49588 9716
rect 49420 9662 49534 9714
rect 49586 9662 49588 9714
rect 49420 9660 49588 9662
rect 49532 9650 49588 9660
rect 49756 9044 49812 9772
rect 49868 9716 49924 9726
rect 49868 9622 49924 9660
rect 49756 8146 49812 8988
rect 49756 8094 49758 8146
rect 49810 8094 49812 8146
rect 49756 8082 49812 8094
rect 49420 7364 49476 7374
rect 49420 7362 49812 7364
rect 49420 7310 49422 7362
rect 49474 7310 49812 7362
rect 49420 7308 49812 7310
rect 49420 7298 49476 7308
rect 49308 7084 49700 7140
rect 49196 7028 49252 7038
rect 48692 6636 48916 6692
rect 48636 6598 48692 6636
rect 48188 6524 48356 6580
rect 48300 6468 48356 6524
rect 48636 6468 48692 6478
rect 48300 6466 48692 6468
rect 48300 6414 48638 6466
rect 48690 6414 48692 6466
rect 48300 6412 48692 6414
rect 47852 6402 47908 6412
rect 48636 6402 48692 6412
rect 48748 5906 48804 6636
rect 48860 6578 48916 6636
rect 48860 6526 48862 6578
rect 48914 6526 48916 6578
rect 48860 6514 48916 6526
rect 48748 5854 48750 5906
rect 48802 5854 48804 5906
rect 48748 5842 48804 5854
rect 49196 5908 49252 6972
rect 49532 6580 49588 6590
rect 49532 6486 49588 6524
rect 49196 5906 49588 5908
rect 49196 5854 49198 5906
rect 49250 5854 49588 5906
rect 49196 5852 49588 5854
rect 49196 5842 49252 5852
rect 49532 5234 49588 5852
rect 49532 5182 49534 5234
rect 49586 5182 49588 5234
rect 49532 5170 49588 5182
rect 48860 5124 48916 5134
rect 48860 4562 48916 5068
rect 48860 4510 48862 4562
rect 48914 4510 48916 4562
rect 48860 4498 48916 4510
rect 49420 4564 49476 4574
rect 49644 4564 49700 7084
rect 49756 6690 49812 7308
rect 49980 6914 50036 9884
rect 50204 9716 50260 9726
rect 50092 9714 50260 9716
rect 50092 9662 50206 9714
rect 50258 9662 50260 9714
rect 50092 9660 50260 9662
rect 50092 9604 50148 9660
rect 50204 9650 50260 9660
rect 50092 7474 50148 9548
rect 50092 7422 50094 7474
rect 50146 7422 50148 7474
rect 50092 7410 50148 7422
rect 50204 7588 50260 7598
rect 50204 7362 50260 7532
rect 50204 7310 50206 7362
rect 50258 7310 50260 7362
rect 50204 7298 50260 7310
rect 49980 6862 49982 6914
rect 50034 6862 50036 6914
rect 49980 6804 50036 6862
rect 49980 6738 50036 6748
rect 49756 6638 49758 6690
rect 49810 6638 49812 6690
rect 49756 6626 49812 6638
rect 50204 6690 50260 6702
rect 50204 6638 50206 6690
rect 50258 6638 50260 6690
rect 50204 6468 50260 6638
rect 50204 6402 50260 6412
rect 50316 5906 50372 10556
rect 50540 9716 50596 9726
rect 50540 9622 50596 9660
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50428 7588 50484 7598
rect 50428 6690 50484 7532
rect 50428 6638 50430 6690
rect 50482 6638 50484 6690
rect 50428 6626 50484 6638
rect 51548 6692 51604 16604
rect 51884 16098 51940 17052
rect 51884 16046 51886 16098
rect 51938 16046 51940 16098
rect 51884 16034 51940 16046
rect 51772 15876 51828 15886
rect 51772 15426 51828 15820
rect 51772 15374 51774 15426
rect 51826 15374 51828 15426
rect 51772 15362 51828 15374
rect 51996 15876 52052 15886
rect 52108 15876 52164 17948
rect 52556 17444 52612 18398
rect 52780 17556 52836 18956
rect 52892 18946 52948 18956
rect 52780 17490 52836 17500
rect 52892 18450 52948 18462
rect 52892 18398 52894 18450
rect 52946 18398 52948 18450
rect 52556 17378 52612 17388
rect 52892 17220 52948 18398
rect 53004 17668 53060 21644
rect 53228 21606 53284 21644
rect 53228 19908 53284 19918
rect 53228 19814 53284 19852
rect 53228 19348 53284 19358
rect 53228 19234 53284 19292
rect 53228 19182 53230 19234
rect 53282 19182 53284 19234
rect 53228 19170 53284 19182
rect 53004 17602 53060 17612
rect 52892 17164 53060 17220
rect 52892 16996 52948 17006
rect 52892 16902 52948 16940
rect 52668 16884 52724 16894
rect 52668 16790 52724 16828
rect 52556 16156 52948 16212
rect 52220 16100 52276 16110
rect 52556 16100 52612 16156
rect 52220 16098 52612 16100
rect 52220 16046 52222 16098
rect 52274 16046 52612 16098
rect 52220 16044 52612 16046
rect 52892 16098 52948 16156
rect 52892 16046 52894 16098
rect 52946 16046 52948 16098
rect 52220 16034 52276 16044
rect 52892 16034 52948 16046
rect 53004 16100 53060 17164
rect 53228 16884 53284 16894
rect 53228 16790 53284 16828
rect 53116 16100 53172 16110
rect 53004 16098 53172 16100
rect 53004 16046 53118 16098
rect 53170 16046 53172 16098
rect 53004 16044 53172 16046
rect 52668 15988 52724 15998
rect 52668 15894 52724 15932
rect 51996 15874 52164 15876
rect 51996 15822 51998 15874
rect 52050 15822 52164 15874
rect 51996 15820 52164 15822
rect 52780 15876 52836 15886
rect 51996 12068 52052 15820
rect 52780 15782 52836 15820
rect 52332 15540 52388 15550
rect 52332 15446 52388 15484
rect 53116 15428 53172 16044
rect 53116 15362 53172 15372
rect 52108 15204 52164 15242
rect 52108 15138 52164 15148
rect 52220 15202 52276 15214
rect 52220 15150 52222 15202
rect 52274 15150 52276 15202
rect 52220 13524 52276 15150
rect 52668 15092 52724 15102
rect 52668 14642 52724 15036
rect 52668 14590 52670 14642
rect 52722 14590 52724 14642
rect 52668 14578 52724 14590
rect 52220 13458 52276 13468
rect 52668 14420 52724 14430
rect 51996 12002 52052 12012
rect 52220 11284 52276 11294
rect 52220 11190 52276 11228
rect 52220 9044 52276 9054
rect 52220 8950 52276 8988
rect 52556 8818 52612 8830
rect 52556 8766 52558 8818
rect 52610 8766 52612 8818
rect 52332 7588 52388 7598
rect 52332 7494 52388 7532
rect 52556 7476 52612 8766
rect 52668 8428 52724 14364
rect 52892 14308 52948 14318
rect 52892 11282 52948 14252
rect 53228 14306 53284 14318
rect 53228 14254 53230 14306
rect 53282 14254 53284 14306
rect 53228 13972 53284 14254
rect 53340 13972 53396 13982
rect 53228 13916 53340 13972
rect 53340 13878 53396 13916
rect 53228 12068 53284 12078
rect 53228 11974 53284 12012
rect 52892 11230 52894 11282
rect 52946 11230 52948 11282
rect 52892 11218 52948 11230
rect 53228 11284 53284 11294
rect 53228 11190 53284 11228
rect 53228 10500 53284 10510
rect 52780 10498 53284 10500
rect 52780 10446 53230 10498
rect 53282 10446 53284 10498
rect 52780 10444 53284 10446
rect 52780 9716 52836 10444
rect 53228 10434 53284 10444
rect 52780 9042 52836 9660
rect 52780 8990 52782 9042
rect 52834 8990 52836 9042
rect 52780 8978 52836 8990
rect 53228 8596 53284 8606
rect 52668 8372 52948 8428
rect 52892 8146 52948 8372
rect 53228 8260 53284 8540
rect 53228 8258 53396 8260
rect 53228 8206 53230 8258
rect 53282 8206 53396 8258
rect 53228 8204 53396 8206
rect 53228 8194 53284 8204
rect 52892 8094 52894 8146
rect 52946 8094 52948 8146
rect 52892 8082 52948 8094
rect 53340 7698 53396 8204
rect 53340 7646 53342 7698
rect 53394 7646 53396 7698
rect 53340 7634 53396 7646
rect 52668 7476 52724 7486
rect 52556 7474 52836 7476
rect 52556 7422 52670 7474
rect 52722 7422 52836 7474
rect 52556 7420 52836 7422
rect 52668 7410 52724 7420
rect 51548 6626 51604 6636
rect 52668 6692 52724 6702
rect 52668 6598 52724 6636
rect 50764 6580 50820 6590
rect 50540 6578 50820 6580
rect 50540 6526 50766 6578
rect 50818 6526 50820 6578
rect 50540 6524 50820 6526
rect 50540 6466 50596 6524
rect 50764 6514 50820 6524
rect 50540 6414 50542 6466
rect 50594 6414 50596 6466
rect 50540 6402 50596 6414
rect 50876 6468 50932 6478
rect 52220 6468 52276 6478
rect 50876 6466 51156 6468
rect 50876 6414 50878 6466
rect 50930 6414 51156 6466
rect 50876 6412 51156 6414
rect 50876 6402 50932 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 51100 6018 51156 6412
rect 52220 6374 52276 6412
rect 51100 5966 51102 6018
rect 51154 5966 51156 6018
rect 51100 5954 51156 5966
rect 50316 5854 50318 5906
rect 50370 5854 50372 5906
rect 49980 5794 50036 5806
rect 49980 5742 49982 5794
rect 50034 5742 50036 5794
rect 49980 5124 50036 5742
rect 50316 5124 50372 5854
rect 52780 5796 52836 7420
rect 53228 6468 53284 6478
rect 53284 6412 53396 6468
rect 53228 6374 53284 6412
rect 53340 5908 53396 6412
rect 53340 5842 53396 5852
rect 53228 5796 53284 5806
rect 52780 5794 53284 5796
rect 52780 5742 53230 5794
rect 53282 5742 53284 5794
rect 52780 5740 53284 5742
rect 53228 5730 53284 5740
rect 50036 5068 50372 5124
rect 49980 5030 50036 5068
rect 49420 4562 49700 4564
rect 49420 4510 49422 4562
rect 49474 4510 49700 4562
rect 49420 4508 49700 4510
rect 49420 4498 49476 4508
rect 47628 4398 47630 4450
rect 47682 4398 47684 4450
rect 47628 4386 47684 4398
rect 49644 4450 49700 4508
rect 49644 4398 49646 4450
rect 49698 4398 49700 4450
rect 49644 4386 49700 4398
rect 49980 4452 50036 4462
rect 49980 4358 50036 4396
rect 50316 4338 50372 5068
rect 52668 5012 52724 5022
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 51100 4452 51156 4462
rect 51100 4358 51156 4396
rect 50316 4286 50318 4338
rect 50370 4286 50372 4338
rect 50316 4274 50372 4286
rect 48076 4228 48132 4238
rect 46508 3614 46510 3666
rect 46562 3614 46564 3666
rect 46508 3602 46564 3614
rect 47740 4226 48132 4228
rect 47740 4174 48078 4226
rect 48130 4174 48132 4226
rect 47740 4172 48132 4174
rect 47740 3554 47796 4172
rect 48076 4162 48132 4172
rect 50652 3892 50708 3902
rect 49644 3668 49700 3678
rect 49644 3574 49700 3612
rect 47740 3502 47742 3554
rect 47794 3502 47796 3554
rect 44156 3378 44212 3388
rect 47404 3444 47460 3482
rect 47740 3388 47796 3502
rect 50652 3554 50708 3836
rect 50652 3502 50654 3554
rect 50706 3502 50708 3554
rect 50652 3490 50708 3502
rect 51996 3668 52052 3678
rect 47404 3378 47460 3388
rect 42812 2212 42868 3332
rect 47516 3332 47796 3388
rect 42812 2156 43092 2212
rect 43036 800 43092 2156
rect 47516 800 47572 3332
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51996 800 52052 3612
rect 52668 3666 52724 4956
rect 53228 4226 53284 4238
rect 53228 4174 53230 4226
rect 53282 4174 53284 4226
rect 53228 3892 53284 4174
rect 53228 3826 53284 3836
rect 52668 3614 52670 3666
rect 52722 3614 52724 3666
rect 52668 3602 52724 3614
rect 52444 3442 52500 3454
rect 52444 3390 52446 3442
rect 52498 3390 52500 3442
rect 52444 3220 52500 3390
rect 52444 3154 52500 3164
rect 53228 3442 53284 3454
rect 53228 3390 53230 3442
rect 53282 3390 53284 3442
rect 53228 3220 53284 3390
rect 53228 3154 53284 3164
rect 2688 0 2800 800
rect 7168 0 7280 800
rect 11648 0 11760 800
rect 16128 0 16240 800
rect 20608 0 20720 800
rect 25088 0 25200 800
rect 29568 0 29680 800
rect 34048 0 34160 800
rect 38528 0 38640 800
rect 43008 0 43120 800
rect 47488 0 47600 800
rect 51968 0 52080 800
<< via2 >>
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51100 51548 51156 51604
rect 49868 51324 49924 51380
rect 16940 50594 16996 50596
rect 16940 50542 16942 50594
rect 16942 50542 16994 50594
rect 16994 50542 16996 50594
rect 16940 50540 16996 50542
rect 17948 50540 18004 50596
rect 17612 50482 17668 50484
rect 17612 50430 17614 50482
rect 17614 50430 17666 50482
rect 17666 50430 17668 50482
rect 17612 50428 17668 50430
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 7308 45388 7364 45444
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 10444 45778 10500 45780
rect 10444 45726 10446 45778
rect 10446 45726 10498 45778
rect 10498 45726 10500 45778
rect 10444 45724 10500 45726
rect 9772 45388 9828 45444
rect 9660 44434 9716 44436
rect 9660 44382 9662 44434
rect 9662 44382 9714 44434
rect 9714 44382 9716 44434
rect 9660 44380 9716 44382
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 7532 43596 7588 43652
rect 9660 44044 9716 44100
rect 9996 43820 10052 43876
rect 9772 43650 9828 43652
rect 9772 43598 9774 43650
rect 9774 43598 9826 43650
rect 9826 43598 9828 43650
rect 9772 43596 9828 43598
rect 11228 45724 11284 45780
rect 11116 45276 11172 45332
rect 12348 45276 12404 45332
rect 12236 45218 12292 45220
rect 12236 45166 12238 45218
rect 12238 45166 12290 45218
rect 12290 45166 12292 45218
rect 12236 45164 12292 45166
rect 10892 44492 10948 44548
rect 10444 44380 10500 44436
rect 10780 44098 10836 44100
rect 10780 44046 10782 44098
rect 10782 44046 10834 44098
rect 10834 44046 10836 44098
rect 10780 44044 10836 44046
rect 11564 44940 11620 44996
rect 11340 44322 11396 44324
rect 11340 44270 11342 44322
rect 11342 44270 11394 44322
rect 11394 44270 11396 44322
rect 11340 44268 11396 44270
rect 10892 43932 10948 43988
rect 11788 44492 11844 44548
rect 11900 44380 11956 44436
rect 11452 43820 11508 43876
rect 12460 45106 12516 45108
rect 12460 45054 12462 45106
rect 12462 45054 12514 45106
rect 12514 45054 12516 45106
rect 12460 45052 12516 45054
rect 13020 47404 13076 47460
rect 13692 46562 13748 46564
rect 13692 46510 13694 46562
rect 13694 46510 13746 46562
rect 13746 46510 13748 46562
rect 13692 46508 13748 46510
rect 12572 44940 12628 44996
rect 12684 45164 12740 45220
rect 12572 44380 12628 44436
rect 12908 45218 12964 45220
rect 12908 45166 12910 45218
rect 12910 45166 12962 45218
rect 12962 45166 12964 45218
rect 12908 45164 12964 45166
rect 12684 44322 12740 44324
rect 12684 44270 12686 44322
rect 12686 44270 12738 44322
rect 12738 44270 12740 44322
rect 12684 44268 12740 44270
rect 12796 44828 12852 44884
rect 12908 44492 12964 44548
rect 13356 44380 13412 44436
rect 12796 44156 12852 44212
rect 13580 44156 13636 44212
rect 12012 43820 12068 43876
rect 10892 43538 10948 43540
rect 10892 43486 10894 43538
rect 10894 43486 10946 43538
rect 10946 43486 10948 43538
rect 10892 43484 10948 43486
rect 11788 43484 11844 43540
rect 11676 42194 11732 42196
rect 11676 42142 11678 42194
rect 11678 42142 11730 42194
rect 11730 42142 11732 42194
rect 11676 42140 11732 42142
rect 8092 41804 8148 41860
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5740 39618 5796 39620
rect 5740 39566 5742 39618
rect 5742 39566 5794 39618
rect 5794 39566 5796 39618
rect 5740 39564 5796 39566
rect 10220 41132 10276 41188
rect 7308 39564 7364 39620
rect 6524 38834 6580 38836
rect 6524 38782 6526 38834
rect 6526 38782 6578 38834
rect 6578 38782 6580 38834
rect 6524 38780 6580 38782
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2492 37154 2548 37156
rect 2492 37102 2494 37154
rect 2494 37102 2546 37154
rect 2546 37102 2548 37154
rect 2492 37100 2548 37102
rect 5292 37266 5348 37268
rect 5292 37214 5294 37266
rect 5294 37214 5346 37266
rect 5346 37214 5348 37266
rect 5292 37212 5348 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1820 34972 1876 35028
rect 2492 34802 2548 34804
rect 2492 34750 2494 34802
rect 2494 34750 2546 34802
rect 2546 34750 2548 34802
rect 2492 34748 2548 34750
rect 5740 37154 5796 37156
rect 5740 37102 5742 37154
rect 5742 37102 5794 37154
rect 5794 37102 5796 37154
rect 5740 37100 5796 37102
rect 5740 35922 5796 35924
rect 5740 35870 5742 35922
rect 5742 35870 5794 35922
rect 5794 35870 5796 35922
rect 5740 35868 5796 35870
rect 5068 35644 5124 35700
rect 6300 36204 6356 36260
rect 4844 34972 4900 35028
rect 5180 35026 5236 35028
rect 5180 34974 5182 35026
rect 5182 34974 5234 35026
rect 5234 34974 5236 35026
rect 5180 34972 5236 34974
rect 4620 34076 4676 34132
rect 5292 34130 5348 34132
rect 5292 34078 5294 34130
rect 5294 34078 5346 34130
rect 5346 34078 5348 34130
rect 5292 34076 5348 34078
rect 6860 37826 6916 37828
rect 6860 37774 6862 37826
rect 6862 37774 6914 37826
rect 6914 37774 6916 37826
rect 6860 37772 6916 37774
rect 7532 37772 7588 37828
rect 6748 37212 6804 37268
rect 6860 37100 6916 37156
rect 7532 37154 7588 37156
rect 7532 37102 7534 37154
rect 7534 37102 7586 37154
rect 7586 37102 7588 37154
rect 7532 37100 7588 37102
rect 8540 37100 8596 37156
rect 8988 39730 9044 39732
rect 8988 39678 8990 39730
rect 8990 39678 9042 39730
rect 9042 39678 9044 39730
rect 8988 39676 9044 39678
rect 10444 41970 10500 41972
rect 10444 41918 10446 41970
rect 10446 41918 10498 41970
rect 10498 41918 10500 41970
rect 10444 41916 10500 41918
rect 10556 41858 10612 41860
rect 10556 41806 10558 41858
rect 10558 41806 10610 41858
rect 10610 41806 10612 41858
rect 10556 41804 10612 41806
rect 10892 41186 10948 41188
rect 10892 41134 10894 41186
rect 10894 41134 10946 41186
rect 10946 41134 10948 41186
rect 10892 41132 10948 41134
rect 10780 40626 10836 40628
rect 10780 40574 10782 40626
rect 10782 40574 10834 40626
rect 10834 40574 10836 40626
rect 10780 40572 10836 40574
rect 11116 41074 11172 41076
rect 11116 41022 11118 41074
rect 11118 41022 11170 41074
rect 11170 41022 11172 41074
rect 11116 41020 11172 41022
rect 10892 40348 10948 40404
rect 11228 40572 11284 40628
rect 10108 39452 10164 39508
rect 9772 38946 9828 38948
rect 9772 38894 9774 38946
rect 9774 38894 9826 38946
rect 9826 38894 9828 38946
rect 9772 38892 9828 38894
rect 11564 39676 11620 39732
rect 11228 39506 11284 39508
rect 11228 39454 11230 39506
rect 11230 39454 11282 39506
rect 11282 39454 11284 39506
rect 11228 39452 11284 39454
rect 11004 39004 11060 39060
rect 9884 37100 9940 37156
rect 6636 35868 6692 35924
rect 6524 35698 6580 35700
rect 6524 35646 6526 35698
rect 6526 35646 6578 35698
rect 6578 35646 6580 35698
rect 6524 35644 6580 35646
rect 6188 34412 6244 34468
rect 6524 34748 6580 34804
rect 6748 34242 6804 34244
rect 6748 34190 6750 34242
rect 6750 34190 6802 34242
rect 6802 34190 6804 34242
rect 6748 34188 6804 34190
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4956 32508 5012 32564
rect 1820 32396 1876 32452
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2492 31836 2548 31892
rect 4732 31666 4788 31668
rect 4732 31614 4734 31666
rect 4734 31614 4786 31666
rect 4786 31614 4788 31666
rect 4732 31612 4788 31614
rect 5180 32450 5236 32452
rect 5180 32398 5182 32450
rect 5182 32398 5234 32450
rect 5234 32398 5236 32450
rect 5180 32396 5236 32398
rect 5068 31500 5124 31556
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4620 30322 4676 30324
rect 4620 30270 4622 30322
rect 4622 30270 4674 30322
rect 4674 30270 4676 30322
rect 4620 30268 4676 30270
rect 6972 33628 7028 33684
rect 5740 33404 5796 33460
rect 5628 32562 5684 32564
rect 5628 32510 5630 32562
rect 5630 32510 5682 32562
rect 5682 32510 5684 32562
rect 5628 32508 5684 32510
rect 5292 31612 5348 31668
rect 5852 31890 5908 31892
rect 5852 31838 5854 31890
rect 5854 31838 5906 31890
rect 5906 31838 5908 31890
rect 5852 31836 5908 31838
rect 2492 30098 2548 30100
rect 2492 30046 2494 30098
rect 2494 30046 2546 30098
rect 2546 30046 2548 30098
rect 2492 30044 2548 30046
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4956 27858 5012 27860
rect 4956 27806 4958 27858
rect 4958 27806 5010 27858
rect 5010 27806 5012 27858
rect 4956 27804 5012 27806
rect 2492 27746 2548 27748
rect 2492 27694 2494 27746
rect 2494 27694 2546 27746
rect 2546 27694 2548 27746
rect 2492 27692 2548 27694
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 6412 32450 6468 32452
rect 6412 32398 6414 32450
rect 6414 32398 6466 32450
rect 6466 32398 6468 32450
rect 6412 32396 6468 32398
rect 6300 31836 6356 31892
rect 6748 31554 6804 31556
rect 6748 31502 6750 31554
rect 6750 31502 6802 31554
rect 6802 31502 6804 31554
rect 6748 31500 6804 31502
rect 5628 30940 5684 30996
rect 6300 30940 6356 30996
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 2940 25228 2996 25284
rect 5740 30268 5796 30324
rect 5740 28642 5796 28644
rect 5740 28590 5742 28642
rect 5742 28590 5794 28642
rect 5794 28590 5796 28642
rect 5740 28588 5796 28590
rect 5292 28028 5348 28084
rect 5964 28028 6020 28084
rect 6300 30098 6356 30100
rect 6300 30046 6302 30098
rect 6302 30046 6354 30098
rect 6354 30046 6356 30098
rect 6300 30044 6356 30046
rect 6412 29426 6468 29428
rect 6412 29374 6414 29426
rect 6414 29374 6466 29426
rect 6466 29374 6468 29426
rect 6412 29372 6468 29374
rect 6972 30156 7028 30212
rect 6748 30098 6804 30100
rect 6748 30046 6750 30098
rect 6750 30046 6802 30098
rect 6802 30046 6804 30098
rect 6748 30044 6804 30046
rect 6860 29650 6916 29652
rect 6860 29598 6862 29650
rect 6862 29598 6914 29650
rect 6914 29598 6916 29650
rect 6860 29596 6916 29598
rect 6748 29426 6804 29428
rect 6748 29374 6750 29426
rect 6750 29374 6802 29426
rect 6802 29374 6804 29426
rect 6748 29372 6804 29374
rect 7196 34242 7252 34244
rect 7196 34190 7198 34242
rect 7198 34190 7250 34242
rect 7250 34190 7252 34242
rect 7196 34188 7252 34190
rect 8428 35026 8484 35028
rect 8428 34974 8430 35026
rect 8430 34974 8482 35026
rect 8482 34974 8484 35026
rect 8428 34972 8484 34974
rect 9548 36876 9604 36932
rect 8988 34972 9044 35028
rect 9212 36258 9268 36260
rect 9212 36206 9214 36258
rect 9214 36206 9266 36258
rect 9266 36206 9268 36258
rect 9212 36204 9268 36206
rect 9548 35810 9604 35812
rect 9548 35758 9550 35810
rect 9550 35758 9602 35810
rect 9602 35758 9604 35810
rect 9548 35756 9604 35758
rect 9996 36258 10052 36260
rect 9996 36206 9998 36258
rect 9998 36206 10050 36258
rect 10050 36206 10052 36258
rect 9996 36204 10052 36206
rect 9996 35922 10052 35924
rect 9996 35870 9998 35922
rect 9998 35870 10050 35922
rect 10050 35870 10052 35922
rect 9996 35868 10052 35870
rect 9772 35698 9828 35700
rect 9772 35646 9774 35698
rect 9774 35646 9826 35698
rect 9826 35646 9828 35698
rect 9772 35644 9828 35646
rect 9212 34860 9268 34916
rect 7532 34636 7588 34692
rect 8092 34412 8148 34468
rect 7532 34300 7588 34356
rect 7868 34300 7924 34356
rect 7420 34076 7476 34132
rect 7532 31836 7588 31892
rect 7980 33458 8036 33460
rect 7980 33406 7982 33458
rect 7982 33406 8034 33458
rect 8034 33406 8036 33458
rect 7980 33404 8036 33406
rect 8988 34130 9044 34132
rect 8988 34078 8990 34130
rect 8990 34078 9042 34130
rect 9042 34078 9044 34130
rect 8988 34076 9044 34078
rect 8876 33516 8932 33572
rect 8988 33740 9044 33796
rect 7196 30322 7252 30324
rect 7196 30270 7198 30322
rect 7198 30270 7250 30322
rect 7250 30270 7252 30322
rect 7196 30268 7252 30270
rect 7084 29708 7140 29764
rect 6412 28476 6468 28532
rect 6188 28082 6244 28084
rect 6188 28030 6190 28082
rect 6190 28030 6242 28082
rect 6242 28030 6244 28082
rect 6188 28028 6244 28030
rect 6076 27916 6132 27972
rect 5292 27132 5348 27188
rect 5404 25452 5460 25508
rect 4620 24668 4676 24724
rect 5404 24722 5460 24724
rect 5404 24670 5406 24722
rect 5406 24670 5458 24722
rect 5458 24670 5460 24722
rect 5404 24668 5460 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5628 25506 5684 25508
rect 5628 25454 5630 25506
rect 5630 25454 5682 25506
rect 5682 25454 5684 25506
rect 5628 25452 5684 25454
rect 5852 26460 5908 26516
rect 6076 26236 6132 26292
rect 6636 28028 6692 28084
rect 6524 27580 6580 27636
rect 6636 27298 6692 27300
rect 6636 27246 6638 27298
rect 6638 27246 6690 27298
rect 6690 27246 6692 27298
rect 6636 27244 6692 27246
rect 6524 27186 6580 27188
rect 6524 27134 6526 27186
rect 6526 27134 6578 27186
rect 6578 27134 6580 27186
rect 6524 27132 6580 27134
rect 6636 26514 6692 26516
rect 6636 26462 6638 26514
rect 6638 26462 6690 26514
rect 6690 26462 6692 26514
rect 6636 26460 6692 26462
rect 6524 26290 6580 26292
rect 6524 26238 6526 26290
rect 6526 26238 6578 26290
rect 6578 26238 6580 26290
rect 6524 26236 6580 26238
rect 7196 28476 7252 28532
rect 6860 27746 6916 27748
rect 6860 27694 6862 27746
rect 6862 27694 6914 27746
rect 6914 27694 6916 27746
rect 6860 27692 6916 27694
rect 7308 27244 7364 27300
rect 7532 28082 7588 28084
rect 7532 28030 7534 28082
rect 7534 28030 7586 28082
rect 7586 28030 7588 28082
rect 7532 28028 7588 28030
rect 7756 30156 7812 30212
rect 8204 31500 8260 31556
rect 8316 30268 8372 30324
rect 8652 30156 8708 30212
rect 8428 30044 8484 30100
rect 8876 29372 8932 29428
rect 8988 29314 9044 29316
rect 8988 29262 8990 29314
rect 8990 29262 9042 29314
rect 9042 29262 9044 29314
rect 8988 29260 9044 29262
rect 8428 28642 8484 28644
rect 8428 28590 8430 28642
rect 8430 28590 8482 28642
rect 8482 28590 8484 28642
rect 8428 28588 8484 28590
rect 7756 27970 7812 27972
rect 7756 27918 7758 27970
rect 7758 27918 7810 27970
rect 7810 27918 7812 27970
rect 7756 27916 7812 27918
rect 8540 27804 8596 27860
rect 8316 27580 8372 27636
rect 6076 25564 6132 25620
rect 5964 25282 6020 25284
rect 5964 25230 5966 25282
rect 5966 25230 6018 25282
rect 6018 25230 6020 25282
rect 5964 25228 6020 25230
rect 2716 23714 2772 23716
rect 2716 23662 2718 23714
rect 2718 23662 2770 23714
rect 2770 23662 2772 23714
rect 2716 23660 2772 23662
rect 3388 23660 3444 23716
rect 2940 22092 2996 22148
rect 1708 20188 1764 20244
rect 5964 23714 6020 23716
rect 5964 23662 5966 23714
rect 5966 23662 6018 23714
rect 6018 23662 6020 23714
rect 5964 23660 6020 23662
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 6972 26236 7028 26292
rect 6636 23660 6692 23716
rect 7196 23436 7252 23492
rect 9660 34636 9716 34692
rect 10668 36258 10724 36260
rect 10668 36206 10670 36258
rect 10670 36206 10722 36258
rect 10722 36206 10724 36258
rect 10668 36204 10724 36206
rect 10668 35420 10724 35476
rect 10332 34914 10388 34916
rect 10332 34862 10334 34914
rect 10334 34862 10386 34914
rect 10386 34862 10388 34914
rect 10332 34860 10388 34862
rect 9660 33906 9716 33908
rect 9660 33854 9662 33906
rect 9662 33854 9714 33906
rect 9714 33854 9716 33906
rect 9660 33852 9716 33854
rect 9548 33740 9604 33796
rect 9660 33628 9716 33684
rect 11004 34690 11060 34692
rect 11004 34638 11006 34690
rect 11006 34638 11058 34690
rect 11058 34638 11060 34690
rect 11004 34636 11060 34638
rect 10444 34300 10500 34356
rect 9772 33516 9828 33572
rect 9436 32396 9492 32452
rect 10220 33068 10276 33124
rect 11004 33068 11060 33124
rect 10892 31836 10948 31892
rect 9884 30940 9940 30996
rect 9548 29372 9604 29428
rect 10220 30994 10276 30996
rect 10220 30942 10222 30994
rect 10222 30942 10274 30994
rect 10274 30942 10276 30994
rect 10220 30940 10276 30942
rect 9884 29260 9940 29316
rect 10444 29260 10500 29316
rect 10780 29426 10836 29428
rect 10780 29374 10782 29426
rect 10782 29374 10834 29426
rect 10834 29374 10836 29426
rect 10780 29372 10836 29374
rect 9660 28700 9716 28756
rect 10220 28754 10276 28756
rect 10220 28702 10222 28754
rect 10222 28702 10274 28754
rect 10274 28702 10276 28754
rect 10220 28700 10276 28702
rect 10668 28476 10724 28532
rect 9324 28028 9380 28084
rect 10892 29314 10948 29316
rect 10892 29262 10894 29314
rect 10894 29262 10946 29314
rect 10946 29262 10948 29314
rect 10892 29260 10948 29262
rect 11004 27244 11060 27300
rect 11004 26796 11060 26852
rect 11004 26012 11060 26068
rect 9324 25564 9380 25620
rect 9436 25452 9492 25508
rect 9548 25340 9604 25396
rect 5180 22316 5236 22372
rect 5292 21980 5348 22036
rect 5404 21810 5460 21812
rect 5404 21758 5406 21810
rect 5406 21758 5458 21810
rect 5458 21758 5460 21810
rect 5404 21756 5460 21758
rect 5852 22258 5908 22260
rect 5852 22206 5854 22258
rect 5854 22206 5906 22258
rect 5906 22206 5908 22258
rect 5852 22204 5908 22206
rect 3052 20524 3108 20580
rect 2828 20130 2884 20132
rect 2828 20078 2830 20130
rect 2830 20078 2882 20130
rect 2882 20078 2884 20130
rect 2828 20076 2884 20078
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4844 20188 4900 20244
rect 3500 20130 3556 20132
rect 3500 20078 3502 20130
rect 3502 20078 3554 20130
rect 3554 20078 3556 20130
rect 3500 20076 3556 20078
rect 4956 19964 5012 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5180 20018 5236 20020
rect 5180 19966 5182 20018
rect 5182 19966 5234 20018
rect 5234 19966 5236 20018
rect 5180 19964 5236 19966
rect 5964 22146 6020 22148
rect 5964 22094 5966 22146
rect 5966 22094 6018 22146
rect 6018 22094 6020 22146
rect 5964 22092 6020 22094
rect 6076 21980 6132 22036
rect 5852 21698 5908 21700
rect 5852 21646 5854 21698
rect 5854 21646 5906 21698
rect 5906 21646 5908 21698
rect 5852 21644 5908 21646
rect 6188 21644 6244 21700
rect 7532 22988 7588 23044
rect 7084 22316 7140 22372
rect 6636 21586 6692 21588
rect 6636 21534 6638 21586
rect 6638 21534 6690 21586
rect 6690 21534 6692 21586
rect 6636 21532 6692 21534
rect 6300 21474 6356 21476
rect 6300 21422 6302 21474
rect 6302 21422 6354 21474
rect 6354 21422 6356 21474
rect 6300 21420 6356 21422
rect 7644 22316 7700 22372
rect 7308 21698 7364 21700
rect 7308 21646 7310 21698
rect 7310 21646 7362 21698
rect 7362 21646 7364 21698
rect 7308 21644 7364 21646
rect 7756 22258 7812 22260
rect 7756 22206 7758 22258
rect 7758 22206 7810 22258
rect 7810 22206 7812 22258
rect 7756 22204 7812 22206
rect 8092 23436 8148 23492
rect 8316 22594 8372 22596
rect 8316 22542 8318 22594
rect 8318 22542 8370 22594
rect 8370 22542 8372 22594
rect 8316 22540 8372 22542
rect 9660 25564 9716 25620
rect 10332 25394 10388 25396
rect 10332 25342 10334 25394
rect 10334 25342 10386 25394
rect 10386 25342 10388 25394
rect 10332 25340 10388 25342
rect 10668 25394 10724 25396
rect 10668 25342 10670 25394
rect 10670 25342 10722 25394
rect 10722 25342 10724 25394
rect 10668 25340 10724 25342
rect 11676 39004 11732 39060
rect 12236 42028 12292 42084
rect 12124 41020 12180 41076
rect 13020 42082 13076 42084
rect 13020 42030 13022 42082
rect 13022 42030 13074 42082
rect 13074 42030 13076 42082
rect 13020 42028 13076 42030
rect 12908 41970 12964 41972
rect 12908 41918 12910 41970
rect 12910 41918 12962 41970
rect 12962 41918 12964 41970
rect 12908 41916 12964 41918
rect 12684 41186 12740 41188
rect 12684 41134 12686 41186
rect 12686 41134 12738 41186
rect 12738 41134 12740 41186
rect 12684 41132 12740 41134
rect 12572 41020 12628 41076
rect 12908 41074 12964 41076
rect 12908 41022 12910 41074
rect 12910 41022 12962 41074
rect 12962 41022 12964 41074
rect 12908 41020 12964 41022
rect 11788 36876 11844 36932
rect 11900 40348 11956 40404
rect 11788 35868 11844 35924
rect 13692 41916 13748 41972
rect 13692 41186 13748 41188
rect 13692 41134 13694 41186
rect 13694 41134 13746 41186
rect 13746 41134 13748 41186
rect 13692 41132 13748 41134
rect 16268 47458 16324 47460
rect 16268 47406 16270 47458
rect 16270 47406 16322 47458
rect 16322 47406 16324 47458
rect 16268 47404 16324 47406
rect 23100 50706 23156 50708
rect 23100 50654 23102 50706
rect 23102 50654 23154 50706
rect 23154 50654 23156 50706
rect 23100 50652 23156 50654
rect 26124 50652 26180 50708
rect 20188 50594 20244 50596
rect 20188 50542 20190 50594
rect 20190 50542 20242 50594
rect 20242 50542 20244 50594
rect 20188 50540 20244 50542
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19628 49980 19684 50036
rect 20412 49980 20468 50036
rect 19852 49868 19908 49924
rect 20076 49586 20132 49588
rect 20076 49534 20078 49586
rect 20078 49534 20130 49586
rect 20130 49534 20132 49586
rect 20076 49532 20132 49534
rect 21420 50482 21476 50484
rect 21420 50430 21422 50482
rect 21422 50430 21474 50482
rect 21474 50430 21476 50482
rect 21420 50428 21476 50430
rect 21196 50034 21252 50036
rect 21196 49982 21198 50034
rect 21198 49982 21250 50034
rect 21250 49982 21252 50034
rect 21196 49980 21252 49982
rect 21308 49810 21364 49812
rect 21308 49758 21310 49810
rect 21310 49758 21362 49810
rect 21362 49758 21364 49810
rect 21308 49756 21364 49758
rect 21868 50482 21924 50484
rect 21868 50430 21870 50482
rect 21870 50430 21922 50482
rect 21922 50430 21924 50482
rect 21868 50428 21924 50430
rect 22092 50428 22148 50484
rect 22988 50482 23044 50484
rect 22988 50430 22990 50482
rect 22990 50430 23042 50482
rect 23042 50430 23044 50482
rect 22988 50428 23044 50430
rect 21644 49532 21700 49588
rect 20748 49026 20804 49028
rect 20748 48974 20750 49026
rect 20750 48974 20802 49026
rect 20802 48974 20804 49026
rect 20748 48972 20804 48974
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 17948 47404 18004 47460
rect 16940 47346 16996 47348
rect 16940 47294 16942 47346
rect 16942 47294 16994 47346
rect 16994 47294 16996 47346
rect 16940 47292 16996 47294
rect 17948 46898 18004 46900
rect 17948 46846 17950 46898
rect 17950 46846 18002 46898
rect 18002 46846 18004 46898
rect 17948 46844 18004 46846
rect 15820 46620 15876 46676
rect 13916 45724 13972 45780
rect 14812 45724 14868 45780
rect 14252 45106 14308 45108
rect 14252 45054 14254 45106
rect 14254 45054 14306 45106
rect 14306 45054 14308 45106
rect 14252 45052 14308 45054
rect 14140 44156 14196 44212
rect 14476 44156 14532 44212
rect 15148 44156 15204 44212
rect 14700 43932 14756 43988
rect 14812 42476 14868 42532
rect 15484 43260 15540 43316
rect 13804 39788 13860 39844
rect 14140 39788 14196 39844
rect 12124 39340 12180 39396
rect 12012 39228 12068 39284
rect 12796 38946 12852 38948
rect 12796 38894 12798 38946
rect 12798 38894 12850 38946
rect 12850 38894 12852 38946
rect 12796 38892 12852 38894
rect 13916 38892 13972 38948
rect 15484 39676 15540 39732
rect 12460 35756 12516 35812
rect 12012 35420 12068 35476
rect 12124 35308 12180 35364
rect 11900 34412 11956 34468
rect 13356 35532 13412 35588
rect 12796 35420 12852 35476
rect 12460 35308 12516 35364
rect 12236 34188 12292 34244
rect 12012 34130 12068 34132
rect 12012 34078 12014 34130
rect 12014 34078 12066 34130
rect 12066 34078 12068 34130
rect 12012 34076 12068 34078
rect 12684 34130 12740 34132
rect 12684 34078 12686 34130
rect 12686 34078 12738 34130
rect 12738 34078 12740 34130
rect 12684 34076 12740 34078
rect 12572 33964 12628 34020
rect 11228 33516 11284 33572
rect 13580 34242 13636 34244
rect 13580 34190 13582 34242
rect 13582 34190 13634 34242
rect 13634 34190 13636 34242
rect 13580 34188 13636 34190
rect 12908 33964 12964 34020
rect 11788 33068 11844 33124
rect 11340 28700 11396 28756
rect 11452 28476 11508 28532
rect 12684 29314 12740 29316
rect 12684 29262 12686 29314
rect 12686 29262 12738 29314
rect 12738 29262 12740 29314
rect 12684 29260 12740 29262
rect 12124 29036 12180 29092
rect 13692 31890 13748 31892
rect 13692 31838 13694 31890
rect 13694 31838 13746 31890
rect 13746 31838 13748 31890
rect 13692 31836 13748 31838
rect 12908 29650 12964 29652
rect 12908 29598 12910 29650
rect 12910 29598 12962 29650
rect 12962 29598 12964 29650
rect 12908 29596 12964 29598
rect 13020 29314 13076 29316
rect 13020 29262 13022 29314
rect 13022 29262 13074 29314
rect 13074 29262 13076 29314
rect 13020 29260 13076 29262
rect 12796 28924 12852 28980
rect 11900 28700 11956 28756
rect 11228 26236 11284 26292
rect 11340 25340 11396 25396
rect 10444 23548 10500 23604
rect 10220 23436 10276 23492
rect 8316 22370 8372 22372
rect 8316 22318 8318 22370
rect 8318 22318 8370 22370
rect 8370 22318 8372 22370
rect 8316 22316 8372 22318
rect 7980 22258 8036 22260
rect 7980 22206 7982 22258
rect 7982 22206 8034 22258
rect 8034 22206 8036 22258
rect 7980 22204 8036 22206
rect 8988 22316 9044 22372
rect 8764 22204 8820 22260
rect 7868 21756 7924 21812
rect 7420 21532 7476 21588
rect 7196 21420 7252 21476
rect 7756 21084 7812 21140
rect 5740 20578 5796 20580
rect 5740 20526 5742 20578
rect 5742 20526 5794 20578
rect 5794 20526 5796 20578
rect 5740 20524 5796 20526
rect 5628 20018 5684 20020
rect 5628 19966 5630 20018
rect 5630 19966 5682 20018
rect 5682 19966 5684 20018
rect 5628 19964 5684 19966
rect 7084 19740 7140 19796
rect 6860 18508 6916 18564
rect 6636 18396 6692 18452
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 2492 17052 2548 17108
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4956 16492 5012 16548
rect 4620 16156 4676 16212
rect 5628 16492 5684 16548
rect 6188 17666 6244 17668
rect 6188 17614 6190 17666
rect 6190 17614 6242 17666
rect 6242 17614 6244 17666
rect 6188 17612 6244 17614
rect 5404 16156 5460 16212
rect 5292 16044 5348 16100
rect 5068 15986 5124 15988
rect 5068 15934 5070 15986
rect 5070 15934 5122 15986
rect 5122 15934 5124 15986
rect 5068 15932 5124 15934
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4956 13746 5012 13748
rect 4956 13694 4958 13746
rect 4958 13694 5010 13746
rect 5010 13694 5012 13746
rect 4956 13692 5012 13694
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2604 12962 2660 12964
rect 2604 12910 2606 12962
rect 2606 12910 2658 12962
rect 2658 12910 2660 12962
rect 2604 12908 2660 12910
rect 2492 12012 2548 12068
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4620 11564 4676 11620
rect 1820 11116 1876 11172
rect 6412 17106 6468 17108
rect 6412 17054 6414 17106
rect 6414 17054 6466 17106
rect 6466 17054 6468 17106
rect 6412 17052 6468 17054
rect 6300 16492 6356 16548
rect 6188 16156 6244 16212
rect 5964 15932 6020 15988
rect 6076 15426 6132 15428
rect 6076 15374 6078 15426
rect 6078 15374 6130 15426
rect 6130 15374 6132 15426
rect 6076 15372 6132 15374
rect 6748 17388 6804 17444
rect 7532 19068 7588 19124
rect 7532 18508 7588 18564
rect 7196 18172 7252 18228
rect 6860 16828 6916 16884
rect 6636 16492 6692 16548
rect 6524 15484 6580 15540
rect 7420 17666 7476 17668
rect 7420 17614 7422 17666
rect 7422 17614 7474 17666
rect 7474 17614 7476 17666
rect 7420 17612 7476 17614
rect 8092 19852 8148 19908
rect 8652 19906 8708 19908
rect 8652 19854 8654 19906
rect 8654 19854 8706 19906
rect 8706 19854 8708 19906
rect 8652 19852 8708 19854
rect 8204 19740 8260 19796
rect 10108 23324 10164 23380
rect 9324 22204 9380 22260
rect 9996 22258 10052 22260
rect 9996 22206 9998 22258
rect 9998 22206 10050 22258
rect 10050 22206 10052 22258
rect 9996 22204 10052 22206
rect 10668 22540 10724 22596
rect 10780 22370 10836 22372
rect 10780 22318 10782 22370
rect 10782 22318 10834 22370
rect 10834 22318 10836 22370
rect 10780 22316 10836 22318
rect 11340 25116 11396 25172
rect 12460 28476 12516 28532
rect 12908 28812 12964 28868
rect 12012 26684 12068 26740
rect 12908 26908 12964 26964
rect 11788 26124 11844 26180
rect 11564 25900 11620 25956
rect 12348 26290 12404 26292
rect 12348 26238 12350 26290
rect 12350 26238 12402 26290
rect 12402 26238 12404 26290
rect 12348 26236 12404 26238
rect 11900 26012 11956 26068
rect 12348 25900 12404 25956
rect 11676 24834 11732 24836
rect 11676 24782 11678 24834
rect 11678 24782 11730 24834
rect 11730 24782 11732 24834
rect 11676 24780 11732 24782
rect 13132 24946 13188 24948
rect 13132 24894 13134 24946
rect 13134 24894 13186 24946
rect 13186 24894 13188 24946
rect 13132 24892 13188 24894
rect 11676 24610 11732 24612
rect 11676 24558 11678 24610
rect 11678 24558 11730 24610
rect 11730 24558 11732 24610
rect 11676 24556 11732 24558
rect 12684 24722 12740 24724
rect 12684 24670 12686 24722
rect 12686 24670 12738 24722
rect 12738 24670 12740 24722
rect 12684 24668 12740 24670
rect 12796 24610 12852 24612
rect 12796 24558 12798 24610
rect 12798 24558 12850 24610
rect 12850 24558 12852 24610
rect 12796 24556 12852 24558
rect 11228 23548 11284 23604
rect 11340 23436 11396 23492
rect 11452 23378 11508 23380
rect 11452 23326 11454 23378
rect 11454 23326 11506 23378
rect 11506 23326 11508 23378
rect 11452 23324 11508 23326
rect 11564 23212 11620 23268
rect 11564 22930 11620 22932
rect 11564 22878 11566 22930
rect 11566 22878 11618 22930
rect 11618 22878 11620 22930
rect 11564 22876 11620 22878
rect 12908 23324 12964 23380
rect 12684 23266 12740 23268
rect 12684 23214 12686 23266
rect 12686 23214 12738 23266
rect 12738 23214 12740 23266
rect 12684 23212 12740 23214
rect 11340 21084 11396 21140
rect 11900 22316 11956 22372
rect 9660 20188 9716 20244
rect 9884 20300 9940 20356
rect 9324 19852 9380 19908
rect 7980 18396 8036 18452
rect 8316 18450 8372 18452
rect 8316 18398 8318 18450
rect 8318 18398 8370 18450
rect 8370 18398 8372 18450
rect 8316 18396 8372 18398
rect 8316 17442 8372 17444
rect 8316 17390 8318 17442
rect 8318 17390 8370 17442
rect 8370 17390 8372 17442
rect 8316 17388 8372 17390
rect 7532 16828 7588 16884
rect 5292 12460 5348 12516
rect 6412 15036 6468 15092
rect 6860 15036 6916 15092
rect 6636 14754 6692 14756
rect 6636 14702 6638 14754
rect 6638 14702 6690 14754
rect 6690 14702 6692 14754
rect 6636 14700 6692 14702
rect 6636 13916 6692 13972
rect 5628 13746 5684 13748
rect 5628 13694 5630 13746
rect 5630 13694 5682 13746
rect 5682 13694 5684 13746
rect 5628 13692 5684 13694
rect 5740 12460 5796 12516
rect 5404 11452 5460 11508
rect 7420 13970 7476 13972
rect 7420 13918 7422 13970
rect 7422 13918 7474 13970
rect 7474 13918 7476 13970
rect 7420 13916 7476 13918
rect 7532 13858 7588 13860
rect 7532 13806 7534 13858
rect 7534 13806 7586 13858
rect 7586 13806 7588 13858
rect 7532 13804 7588 13806
rect 6860 13356 6916 13412
rect 8988 18450 9044 18452
rect 8988 18398 8990 18450
rect 8990 18398 9042 18450
rect 9042 18398 9044 18450
rect 8988 18396 9044 18398
rect 9100 17778 9156 17780
rect 9100 17726 9102 17778
rect 9102 17726 9154 17778
rect 9154 17726 9156 17778
rect 9100 17724 9156 17726
rect 8092 15036 8148 15092
rect 8316 14700 8372 14756
rect 8204 14306 8260 14308
rect 8204 14254 8206 14306
rect 8206 14254 8258 14306
rect 8258 14254 8260 14306
rect 8204 14252 8260 14254
rect 8092 13692 8148 13748
rect 7644 13356 7700 13412
rect 8204 12908 8260 12964
rect 8652 15426 8708 15428
rect 8652 15374 8654 15426
rect 8654 15374 8706 15426
rect 8706 15374 8708 15426
rect 8652 15372 8708 15374
rect 9548 19292 9604 19348
rect 11340 20860 11396 20916
rect 10556 20188 10612 20244
rect 10220 19794 10276 19796
rect 10220 19742 10222 19794
rect 10222 19742 10274 19794
rect 10274 19742 10276 19794
rect 10220 19740 10276 19742
rect 9772 18396 9828 18452
rect 9660 17836 9716 17892
rect 10108 17778 10164 17780
rect 10108 17726 10110 17778
rect 10110 17726 10162 17778
rect 10162 17726 10164 17778
rect 10108 17724 10164 17726
rect 10668 17778 10724 17780
rect 10668 17726 10670 17778
rect 10670 17726 10722 17778
rect 10722 17726 10724 17778
rect 10668 17724 10724 17726
rect 9660 17666 9716 17668
rect 9660 17614 9662 17666
rect 9662 17614 9714 17666
rect 9714 17614 9716 17666
rect 9660 17612 9716 17614
rect 9660 16098 9716 16100
rect 9660 16046 9662 16098
rect 9662 16046 9714 16098
rect 9714 16046 9716 16098
rect 9660 16044 9716 16046
rect 10220 15820 10276 15876
rect 8876 14252 8932 14308
rect 8764 14140 8820 14196
rect 8652 13746 8708 13748
rect 8652 13694 8654 13746
rect 8654 13694 8706 13746
rect 8706 13694 8708 13746
rect 8652 13692 8708 13694
rect 8428 12850 8484 12852
rect 8428 12798 8430 12850
rect 8430 12798 8482 12850
rect 8482 12798 8484 12850
rect 8428 12796 8484 12798
rect 7868 12460 7924 12516
rect 6860 12348 6916 12404
rect 8428 12402 8484 12404
rect 8428 12350 8430 12402
rect 8430 12350 8482 12402
rect 8482 12350 8484 12402
rect 8428 12348 8484 12350
rect 7420 12178 7476 12180
rect 7420 12126 7422 12178
rect 7422 12126 7474 12178
rect 7474 12126 7476 12178
rect 7420 12124 7476 12126
rect 6524 12066 6580 12068
rect 6524 12014 6526 12066
rect 6526 12014 6578 12066
rect 6578 12014 6580 12066
rect 6524 12012 6580 12014
rect 10332 15484 10388 15540
rect 9212 14588 9268 14644
rect 9660 14642 9716 14644
rect 9660 14590 9662 14642
rect 9662 14590 9714 14642
rect 9714 14590 9716 14642
rect 9660 14588 9716 14590
rect 10108 14588 10164 14644
rect 9436 14140 9492 14196
rect 10108 14028 10164 14084
rect 9100 12796 9156 12852
rect 9212 13804 9268 13860
rect 8988 12012 9044 12068
rect 6412 11900 6468 11956
rect 7644 11954 7700 11956
rect 7644 11902 7646 11954
rect 7646 11902 7698 11954
rect 7698 11902 7700 11954
rect 7644 11900 7700 11902
rect 6188 11618 6244 11620
rect 6188 11566 6190 11618
rect 6190 11566 6242 11618
rect 6242 11566 6244 11618
rect 6188 11564 6244 11566
rect 6412 11506 6468 11508
rect 6412 11454 6414 11506
rect 6414 11454 6466 11506
rect 6466 11454 6468 11506
rect 6412 11452 6468 11454
rect 5068 11170 5124 11172
rect 5068 11118 5070 11170
rect 5070 11118 5122 11170
rect 5122 11118 5124 11170
rect 5068 11116 5124 11118
rect 4284 10444 4340 10500
rect 2156 10332 2212 10388
rect 6300 11228 6356 11284
rect 7084 10610 7140 10612
rect 7084 10558 7086 10610
rect 7086 10558 7138 10610
rect 7138 10558 7140 10610
rect 7084 10556 7140 10558
rect 6188 10498 6244 10500
rect 6188 10446 6190 10498
rect 6190 10446 6242 10498
rect 6242 10446 6244 10498
rect 6188 10444 6244 10446
rect 5628 10332 5684 10388
rect 6524 10386 6580 10388
rect 6524 10334 6526 10386
rect 6526 10334 6578 10386
rect 6578 10334 6580 10386
rect 6524 10332 6580 10334
rect 7420 10332 7476 10388
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 7420 9212 7476 9268
rect 8092 9548 8148 9604
rect 6076 8876 6132 8932
rect 5404 8204 5460 8260
rect 7420 8258 7476 8260
rect 7420 8206 7422 8258
rect 7422 8206 7474 8258
rect 7474 8206 7476 8258
rect 7420 8204 7476 8206
rect 8428 8204 8484 8260
rect 8428 7420 8484 7476
rect 8204 7362 8260 7364
rect 8204 7310 8206 7362
rect 8206 7310 8258 7362
rect 8258 7310 8260 7362
rect 8204 7308 8260 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 3612 6860 3668 6916
rect 8540 7362 8596 7364
rect 8540 7310 8542 7362
rect 8542 7310 8594 7362
rect 8594 7310 8596 7362
rect 8540 7308 8596 7310
rect 9324 11618 9380 11620
rect 9324 11566 9326 11618
rect 9326 11566 9378 11618
rect 9378 11566 9380 11618
rect 9324 11564 9380 11566
rect 10556 15426 10612 15428
rect 10556 15374 10558 15426
rect 10558 15374 10610 15426
rect 10610 15374 10612 15426
rect 10556 15372 10612 15374
rect 11340 20188 11396 20244
rect 13020 23154 13076 23156
rect 13020 23102 13022 23154
rect 13022 23102 13074 23154
rect 13074 23102 13076 23154
rect 13020 23100 13076 23102
rect 13020 22428 13076 22484
rect 13692 29596 13748 29652
rect 13356 28812 13412 28868
rect 13468 28700 13524 28756
rect 14140 36764 14196 36820
rect 14028 35586 14084 35588
rect 14028 35534 14030 35586
rect 14030 35534 14082 35586
rect 14082 35534 14084 35586
rect 14028 35532 14084 35534
rect 13916 27692 13972 27748
rect 14140 31948 14196 32004
rect 13580 24834 13636 24836
rect 13580 24782 13582 24834
rect 13582 24782 13634 24834
rect 13634 24782 13636 24834
rect 13580 24780 13636 24782
rect 13468 24722 13524 24724
rect 13468 24670 13470 24722
rect 13470 24670 13522 24722
rect 13522 24670 13524 24722
rect 13468 24668 13524 24670
rect 14140 29314 14196 29316
rect 14140 29262 14142 29314
rect 14142 29262 14194 29314
rect 14194 29262 14196 29314
rect 14140 29260 14196 29262
rect 14252 26962 14308 26964
rect 14252 26910 14254 26962
rect 14254 26910 14306 26962
rect 14306 26910 14308 26962
rect 14252 26908 14308 26910
rect 15932 45666 15988 45668
rect 15932 45614 15934 45666
rect 15934 45614 15986 45666
rect 15986 45614 15988 45666
rect 15932 45612 15988 45614
rect 15932 44156 15988 44212
rect 16380 46674 16436 46676
rect 16380 46622 16382 46674
rect 16382 46622 16434 46674
rect 16434 46622 16436 46674
rect 16380 46620 16436 46622
rect 16268 46562 16324 46564
rect 16268 46510 16270 46562
rect 16270 46510 16322 46562
rect 16322 46510 16324 46562
rect 16268 46508 16324 46510
rect 17500 46674 17556 46676
rect 17500 46622 17502 46674
rect 17502 46622 17554 46674
rect 17554 46622 17556 46674
rect 17500 46620 17556 46622
rect 16940 45890 16996 45892
rect 16940 45838 16942 45890
rect 16942 45838 16994 45890
rect 16994 45838 16996 45890
rect 16940 45836 16996 45838
rect 17948 45836 18004 45892
rect 17612 45778 17668 45780
rect 17612 45726 17614 45778
rect 17614 45726 17666 45778
rect 17666 45726 17668 45778
rect 17612 45724 17668 45726
rect 16268 45666 16324 45668
rect 16268 45614 16270 45666
rect 16270 45614 16322 45666
rect 16322 45614 16324 45666
rect 16268 45612 16324 45614
rect 16156 43596 16212 43652
rect 16044 42140 16100 42196
rect 16156 40908 16212 40964
rect 17276 44322 17332 44324
rect 17276 44270 17278 44322
rect 17278 44270 17330 44322
rect 17330 44270 17332 44322
rect 17276 44268 17332 44270
rect 16828 44156 16884 44212
rect 16492 44044 16548 44100
rect 16828 43314 16884 43316
rect 16828 43262 16830 43314
rect 16830 43262 16882 43314
rect 16882 43262 16884 43314
rect 16828 43260 16884 43262
rect 16716 43036 16772 43092
rect 17388 44098 17444 44100
rect 17388 44046 17390 44098
rect 17390 44046 17442 44098
rect 17442 44046 17444 44098
rect 17388 44044 17444 44046
rect 17724 44268 17780 44324
rect 17836 45052 17892 45108
rect 17500 43820 17556 43876
rect 17612 43036 17668 43092
rect 17052 42924 17108 42980
rect 17948 43932 18004 43988
rect 16380 37884 16436 37940
rect 17500 39676 17556 39732
rect 16716 37772 16772 37828
rect 15484 36652 15540 36708
rect 15596 35698 15652 35700
rect 15596 35646 15598 35698
rect 15598 35646 15650 35698
rect 15650 35646 15652 35698
rect 15596 35644 15652 35646
rect 15036 34130 15092 34132
rect 15036 34078 15038 34130
rect 15038 34078 15090 34130
rect 15090 34078 15092 34130
rect 15036 34076 15092 34078
rect 14476 33068 14532 33124
rect 14924 32674 14980 32676
rect 14924 32622 14926 32674
rect 14926 32622 14978 32674
rect 14978 32622 14980 32674
rect 14924 32620 14980 32622
rect 15708 34636 15764 34692
rect 15484 33068 15540 33124
rect 15484 32674 15540 32676
rect 15484 32622 15486 32674
rect 15486 32622 15538 32674
rect 15538 32622 15540 32674
rect 15484 32620 15540 32622
rect 15148 32002 15204 32004
rect 15148 31950 15150 32002
rect 15150 31950 15202 32002
rect 15202 31950 15204 32002
rect 15148 31948 15204 31950
rect 16044 35868 16100 35924
rect 16492 36652 16548 36708
rect 16604 35922 16660 35924
rect 16604 35870 16606 35922
rect 16606 35870 16658 35922
rect 16658 35870 16660 35922
rect 16604 35868 16660 35870
rect 16716 35532 16772 35588
rect 16940 35420 16996 35476
rect 16268 33404 16324 33460
rect 15932 31500 15988 31556
rect 16156 31612 16212 31668
rect 13356 23436 13412 23492
rect 13244 22988 13300 23044
rect 13692 22482 13748 22484
rect 13692 22430 13694 22482
rect 13694 22430 13746 22482
rect 13746 22430 13748 22482
rect 13692 22428 13748 22430
rect 13132 22316 13188 22372
rect 13468 22258 13524 22260
rect 13468 22206 13470 22258
rect 13470 22206 13522 22258
rect 13522 22206 13524 22258
rect 13468 22204 13524 22206
rect 14028 22876 14084 22932
rect 13916 22370 13972 22372
rect 13916 22318 13918 22370
rect 13918 22318 13970 22370
rect 13970 22318 13972 22370
rect 13916 22316 13972 22318
rect 14700 24892 14756 24948
rect 14364 23100 14420 23156
rect 15260 26402 15316 26404
rect 15260 26350 15262 26402
rect 15262 26350 15314 26402
rect 15314 26350 15316 26402
rect 15260 26348 15316 26350
rect 14924 23100 14980 23156
rect 14364 22540 14420 22596
rect 14812 22370 14868 22372
rect 14812 22318 14814 22370
rect 14814 22318 14866 22370
rect 14866 22318 14868 22370
rect 14812 22316 14868 22318
rect 11900 20524 11956 20580
rect 11788 20076 11844 20132
rect 11452 19122 11508 19124
rect 11452 19070 11454 19122
rect 11454 19070 11506 19122
rect 11506 19070 11508 19122
rect 11452 19068 11508 19070
rect 11116 16828 11172 16884
rect 13020 20076 13076 20132
rect 12572 18450 12628 18452
rect 12572 18398 12574 18450
rect 12574 18398 12626 18450
rect 12626 18398 12628 18450
rect 12572 18396 12628 18398
rect 11900 16828 11956 16884
rect 12908 16268 12964 16324
rect 12908 15372 12964 15428
rect 11228 15260 11284 15316
rect 10332 11228 10388 11284
rect 10780 14028 10836 14084
rect 13580 18396 13636 18452
rect 15820 30044 15876 30100
rect 15372 22540 15428 22596
rect 15484 29260 15540 29316
rect 14700 20130 14756 20132
rect 14700 20078 14702 20130
rect 14702 20078 14754 20130
rect 14754 20078 14756 20130
rect 14700 20076 14756 20078
rect 15036 20130 15092 20132
rect 15036 20078 15038 20130
rect 15038 20078 15090 20130
rect 15090 20078 15092 20130
rect 15036 20076 15092 20078
rect 14364 17724 14420 17780
rect 14476 18508 14532 18564
rect 13916 16994 13972 16996
rect 13916 16942 13918 16994
rect 13918 16942 13970 16994
rect 13970 16942 13972 16994
rect 13916 16940 13972 16942
rect 13132 16882 13188 16884
rect 13132 16830 13134 16882
rect 13134 16830 13186 16882
rect 13186 16830 13188 16882
rect 13132 16828 13188 16830
rect 13468 16882 13524 16884
rect 13468 16830 13470 16882
rect 13470 16830 13522 16882
rect 13522 16830 13524 16882
rect 13468 16828 13524 16830
rect 13580 16268 13636 16324
rect 13580 16098 13636 16100
rect 13580 16046 13582 16098
rect 13582 16046 13634 16098
rect 13634 16046 13636 16098
rect 13580 16044 13636 16046
rect 13580 15820 13636 15876
rect 13020 14476 13076 14532
rect 11564 14028 11620 14084
rect 11900 13916 11956 13972
rect 13132 14028 13188 14084
rect 12348 13858 12404 13860
rect 12348 13806 12350 13858
rect 12350 13806 12402 13858
rect 12402 13806 12404 13858
rect 12348 13804 12404 13806
rect 11228 12738 11284 12740
rect 11228 12686 11230 12738
rect 11230 12686 11282 12738
rect 11282 12686 11284 12738
rect 11228 12684 11284 12686
rect 14252 15820 14308 15876
rect 14812 17052 14868 17108
rect 14588 16882 14644 16884
rect 14588 16830 14590 16882
rect 14590 16830 14642 16882
rect 14642 16830 14644 16882
rect 14588 16828 14644 16830
rect 14924 16658 14980 16660
rect 14924 16606 14926 16658
rect 14926 16606 14978 16658
rect 14978 16606 14980 16658
rect 14924 16604 14980 16606
rect 14588 15260 14644 15316
rect 16604 31666 16660 31668
rect 16604 31614 16606 31666
rect 16606 31614 16658 31666
rect 16658 31614 16660 31666
rect 16604 31612 16660 31614
rect 16380 31164 16436 31220
rect 16492 30940 16548 30996
rect 16380 30882 16436 30884
rect 16380 30830 16382 30882
rect 16382 30830 16434 30882
rect 16434 30830 16436 30882
rect 16380 30828 16436 30830
rect 16268 29036 16324 29092
rect 16716 30940 16772 30996
rect 19292 46898 19348 46900
rect 19292 46846 19294 46898
rect 19294 46846 19346 46898
rect 19346 46846 19348 46898
rect 19292 46844 19348 46846
rect 18732 46620 18788 46676
rect 18508 45778 18564 45780
rect 18508 45726 18510 45778
rect 18510 45726 18562 45778
rect 18562 45726 18564 45778
rect 18508 45724 18564 45726
rect 19292 44322 19348 44324
rect 19292 44270 19294 44322
rect 19294 44270 19346 44322
rect 19346 44270 19348 44322
rect 19292 44268 19348 44270
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19628 46732 19684 46788
rect 20524 47458 20580 47460
rect 20524 47406 20526 47458
rect 20526 47406 20578 47458
rect 20578 47406 20580 47458
rect 20524 47404 20580 47406
rect 21420 47346 21476 47348
rect 21420 47294 21422 47346
rect 21422 47294 21474 47346
rect 21474 47294 21476 47346
rect 21420 47292 21476 47294
rect 20524 46786 20580 46788
rect 20524 46734 20526 46786
rect 20526 46734 20578 46786
rect 20578 46734 20580 46786
rect 20524 46732 20580 46734
rect 21084 46786 21140 46788
rect 21084 46734 21086 46786
rect 21086 46734 21138 46786
rect 21138 46734 21140 46786
rect 21084 46732 21140 46734
rect 20636 46674 20692 46676
rect 20636 46622 20638 46674
rect 20638 46622 20690 46674
rect 20690 46622 20692 46674
rect 20636 46620 20692 46622
rect 21756 49026 21812 49028
rect 21756 48974 21758 49026
rect 21758 48974 21810 49026
rect 21810 48974 21812 49026
rect 21756 48972 21812 48974
rect 22428 48914 22484 48916
rect 22428 48862 22430 48914
rect 22430 48862 22482 48914
rect 22482 48862 22484 48914
rect 22428 48860 22484 48862
rect 22316 48748 22372 48804
rect 21868 47346 21924 47348
rect 21868 47294 21870 47346
rect 21870 47294 21922 47346
rect 21922 47294 21924 47346
rect 21868 47292 21924 47294
rect 20300 46060 20356 46116
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19516 45106 19572 45108
rect 19516 45054 19518 45106
rect 19518 45054 19570 45106
rect 19570 45054 19572 45106
rect 19516 45052 19572 45054
rect 19852 44882 19908 44884
rect 19852 44830 19854 44882
rect 19854 44830 19906 44882
rect 19906 44830 19908 44882
rect 19852 44828 19908 44830
rect 19740 44716 19796 44772
rect 20076 45164 20132 45220
rect 19068 43708 19124 43764
rect 18956 43260 19012 43316
rect 18060 42476 18116 42532
rect 17948 41244 18004 41300
rect 18060 41074 18116 41076
rect 18060 41022 18062 41074
rect 18062 41022 18114 41074
rect 18114 41022 18116 41074
rect 18060 41020 18116 41022
rect 17836 40348 17892 40404
rect 17836 39676 17892 39732
rect 19180 42754 19236 42756
rect 19180 42702 19182 42754
rect 19182 42702 19234 42754
rect 19234 42702 19236 42754
rect 19180 42700 19236 42702
rect 18732 41186 18788 41188
rect 18732 41134 18734 41186
rect 18734 41134 18786 41186
rect 18786 41134 18788 41186
rect 18732 41132 18788 41134
rect 18508 41074 18564 41076
rect 18508 41022 18510 41074
rect 18510 41022 18562 41074
rect 18562 41022 18564 41074
rect 18508 41020 18564 41022
rect 18620 40962 18676 40964
rect 18620 40910 18622 40962
rect 18622 40910 18674 40962
rect 18674 40910 18676 40962
rect 18620 40908 18676 40910
rect 18172 39676 18228 39732
rect 18396 40348 18452 40404
rect 18956 41020 19012 41076
rect 19068 40402 19124 40404
rect 19068 40350 19070 40402
rect 19070 40350 19122 40402
rect 19122 40350 19124 40402
rect 19068 40348 19124 40350
rect 18956 39730 19012 39732
rect 18956 39678 18958 39730
rect 18958 39678 19010 39730
rect 19010 39678 19012 39730
rect 18956 39676 19012 39678
rect 18956 39340 19012 39396
rect 18172 37324 18228 37380
rect 17948 37212 18004 37268
rect 17836 36876 17892 36932
rect 18844 37266 18900 37268
rect 18844 37214 18846 37266
rect 18846 37214 18898 37266
rect 18898 37214 18900 37266
rect 18844 37212 18900 37214
rect 17500 35026 17556 35028
rect 17500 34974 17502 35026
rect 17502 34974 17554 35026
rect 17554 34974 17556 35026
rect 17500 34972 17556 34974
rect 18284 37100 18340 37156
rect 18172 36764 18228 36820
rect 17388 33068 17444 33124
rect 18172 34690 18228 34692
rect 18172 34638 18174 34690
rect 18174 34638 18226 34690
rect 18226 34638 18228 34690
rect 18172 34636 18228 34638
rect 16940 30828 16996 30884
rect 17276 30098 17332 30100
rect 17276 30046 17278 30098
rect 17278 30046 17330 30098
rect 17330 30046 17332 30098
rect 17276 30044 17332 30046
rect 17276 29596 17332 29652
rect 16828 29314 16884 29316
rect 16828 29262 16830 29314
rect 16830 29262 16882 29314
rect 16882 29262 16884 29314
rect 16828 29260 16884 29262
rect 16492 28754 16548 28756
rect 16492 28702 16494 28754
rect 16494 28702 16546 28754
rect 16546 28702 16548 28754
rect 16492 28700 16548 28702
rect 16268 28588 16324 28644
rect 17724 31218 17780 31220
rect 17724 31166 17726 31218
rect 17726 31166 17778 31218
rect 17778 31166 17780 31218
rect 17724 31164 17780 31166
rect 17948 33122 18004 33124
rect 17948 33070 17950 33122
rect 17950 33070 18002 33122
rect 18002 33070 18004 33122
rect 17948 33068 18004 33070
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20076 43708 20132 43764
rect 19404 43650 19460 43652
rect 19404 43598 19406 43650
rect 19406 43598 19458 43650
rect 19458 43598 19460 43650
rect 19404 43596 19460 43598
rect 19740 43148 19796 43204
rect 20412 43148 20468 43204
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19628 41132 19684 41188
rect 20412 41692 20468 41748
rect 20524 41132 20580 41188
rect 20636 41244 20692 41300
rect 20188 41074 20244 41076
rect 20188 41022 20190 41074
rect 20190 41022 20242 41074
rect 20242 41022 20244 41074
rect 20188 41020 20244 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20524 40684 20580 40740
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19628 37378 19684 37380
rect 19628 37326 19630 37378
rect 19630 37326 19682 37378
rect 19682 37326 19684 37378
rect 19628 37324 19684 37326
rect 19852 37154 19908 37156
rect 19852 37102 19854 37154
rect 19854 37102 19906 37154
rect 19906 37102 19908 37154
rect 19852 37100 19908 37102
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19740 35698 19796 35700
rect 19740 35646 19742 35698
rect 19742 35646 19794 35698
rect 19794 35646 19796 35698
rect 19740 35644 19796 35646
rect 18620 34412 18676 34468
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21644 46114 21700 46116
rect 21644 46062 21646 46114
rect 21646 46062 21698 46114
rect 21698 46062 21700 46114
rect 21644 46060 21700 46062
rect 21980 45276 22036 45332
rect 22988 49756 23044 49812
rect 23436 50428 23492 50484
rect 23324 49922 23380 49924
rect 23324 49870 23326 49922
rect 23326 49870 23378 49922
rect 23378 49870 23380 49922
rect 23324 49868 23380 49870
rect 23996 50482 24052 50484
rect 23996 50430 23998 50482
rect 23998 50430 24050 50482
rect 24050 50430 24052 50482
rect 23996 50428 24052 50430
rect 22876 48802 22932 48804
rect 22876 48750 22878 48802
rect 22878 48750 22930 48802
rect 22930 48750 22932 48802
rect 22876 48748 22932 48750
rect 22764 47628 22820 47684
rect 22428 47404 22484 47460
rect 22316 45164 22372 45220
rect 21980 44716 22036 44772
rect 22092 44434 22148 44436
rect 22092 44382 22094 44434
rect 22094 44382 22146 44434
rect 22146 44382 22148 44434
rect 22092 44380 22148 44382
rect 22428 44994 22484 44996
rect 22428 44942 22430 44994
rect 22430 44942 22482 44994
rect 22482 44942 22484 44994
rect 22428 44940 22484 44942
rect 22316 44716 22372 44772
rect 23548 48972 23604 49028
rect 23660 49084 23716 49140
rect 23996 48860 24052 48916
rect 23548 48636 23604 48692
rect 23660 48188 23716 48244
rect 22764 46620 22820 46676
rect 23212 46674 23268 46676
rect 23212 46622 23214 46674
rect 23214 46622 23266 46674
rect 23266 46622 23268 46674
rect 23212 46620 23268 46622
rect 26348 50706 26404 50708
rect 26348 50654 26350 50706
rect 26350 50654 26402 50706
rect 26402 50654 26404 50706
rect 26348 50652 26404 50654
rect 24332 50428 24388 50484
rect 26012 50428 26068 50484
rect 25900 49922 25956 49924
rect 25900 49870 25902 49922
rect 25902 49870 25954 49922
rect 25954 49870 25956 49922
rect 25900 49868 25956 49870
rect 25564 49084 25620 49140
rect 31276 50706 31332 50708
rect 31276 50654 31278 50706
rect 31278 50654 31330 50706
rect 31330 50654 31332 50706
rect 31276 50652 31332 50654
rect 29148 50428 29204 50484
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 32396 50594 32452 50596
rect 32396 50542 32398 50594
rect 32398 50542 32450 50594
rect 32450 50542 32452 50594
rect 32396 50540 32452 50542
rect 25788 49026 25844 49028
rect 25788 48974 25790 49026
rect 25790 48974 25842 49026
rect 25842 48974 25844 49026
rect 25788 48972 25844 48974
rect 24556 48914 24612 48916
rect 24556 48862 24558 48914
rect 24558 48862 24610 48914
rect 24610 48862 24612 48914
rect 24556 48860 24612 48862
rect 25340 48914 25396 48916
rect 25340 48862 25342 48914
rect 25342 48862 25394 48914
rect 25394 48862 25396 48914
rect 25340 48860 25396 48862
rect 24108 48748 24164 48804
rect 24444 48748 24500 48804
rect 26348 49196 26404 49252
rect 26796 49810 26852 49812
rect 26796 49758 26798 49810
rect 26798 49758 26850 49810
rect 26850 49758 26852 49810
rect 26796 49756 26852 49758
rect 27356 49922 27412 49924
rect 27356 49870 27358 49922
rect 27358 49870 27410 49922
rect 27410 49870 27412 49922
rect 27356 49868 27412 49870
rect 26572 49698 26628 49700
rect 26572 49646 26574 49698
rect 26574 49646 26626 49698
rect 26626 49646 26628 49698
rect 26572 49644 26628 49646
rect 23100 46060 23156 46116
rect 22988 45836 23044 45892
rect 22652 45164 22708 45220
rect 22988 45276 23044 45332
rect 24780 45836 24836 45892
rect 24108 45778 24164 45780
rect 24108 45726 24110 45778
rect 24110 45726 24162 45778
rect 24162 45726 24164 45778
rect 24108 45724 24164 45726
rect 24668 45724 24724 45780
rect 23548 45612 23604 45668
rect 22876 44492 22932 44548
rect 22652 43596 22708 43652
rect 21308 42700 21364 42756
rect 21532 41916 21588 41972
rect 21308 41692 21364 41748
rect 21196 41074 21252 41076
rect 21196 41022 21198 41074
rect 21198 41022 21250 41074
rect 21250 41022 21252 41074
rect 21196 41020 21252 41022
rect 21532 40684 21588 40740
rect 21756 41804 21812 41860
rect 22764 43148 22820 43204
rect 21980 43036 22036 43092
rect 24444 45666 24500 45668
rect 24444 45614 24446 45666
rect 24446 45614 24498 45666
rect 24498 45614 24500 45666
rect 24444 45612 24500 45614
rect 24668 45330 24724 45332
rect 24668 45278 24670 45330
rect 24670 45278 24722 45330
rect 24722 45278 24724 45330
rect 24668 45276 24724 45278
rect 26684 48748 26740 48804
rect 25900 47346 25956 47348
rect 25900 47294 25902 47346
rect 25902 47294 25954 47346
rect 25954 47294 25956 47346
rect 25900 47292 25956 47294
rect 26124 47180 26180 47236
rect 25900 45890 25956 45892
rect 25900 45838 25902 45890
rect 25902 45838 25954 45890
rect 25954 45838 25956 45890
rect 25900 45836 25956 45838
rect 25340 45612 25396 45668
rect 25676 45106 25732 45108
rect 25676 45054 25678 45106
rect 25678 45054 25730 45106
rect 25730 45054 25732 45106
rect 25676 45052 25732 45054
rect 25116 44940 25172 44996
rect 23996 44828 24052 44884
rect 25788 44940 25844 44996
rect 25900 44546 25956 44548
rect 25900 44494 25902 44546
rect 25902 44494 25954 44546
rect 25954 44494 25956 44546
rect 25900 44492 25956 44494
rect 24108 43596 24164 43652
rect 23660 42754 23716 42756
rect 23660 42702 23662 42754
rect 23662 42702 23714 42754
rect 23714 42702 23716 42754
rect 23660 42700 23716 42702
rect 25452 42866 25508 42868
rect 25452 42814 25454 42866
rect 25454 42814 25506 42866
rect 25506 42814 25508 42866
rect 25452 42812 25508 42814
rect 35756 50594 35812 50596
rect 35756 50542 35758 50594
rect 35758 50542 35810 50594
rect 35810 50542 35812 50594
rect 35756 50540 35812 50542
rect 33180 50482 33236 50484
rect 33180 50430 33182 50482
rect 33182 50430 33234 50482
rect 33234 50430 33236 50482
rect 33180 50428 33236 50430
rect 33964 50428 34020 50484
rect 39900 50594 39956 50596
rect 39900 50542 39902 50594
rect 39902 50542 39954 50594
rect 39954 50542 39956 50594
rect 39900 50540 39956 50542
rect 37660 50428 37716 50484
rect 35084 49980 35140 50036
rect 33852 49922 33908 49924
rect 33852 49870 33854 49922
rect 33854 49870 33906 49922
rect 33906 49870 33908 49922
rect 33852 49868 33908 49870
rect 27692 49810 27748 49812
rect 27692 49758 27694 49810
rect 27694 49758 27746 49810
rect 27746 49758 27748 49810
rect 27692 49756 27748 49758
rect 28028 49532 28084 49588
rect 27132 48914 27188 48916
rect 27132 48862 27134 48914
rect 27134 48862 27186 48914
rect 27186 48862 27188 48914
rect 27132 48860 27188 48862
rect 31388 49698 31444 49700
rect 31388 49646 31390 49698
rect 31390 49646 31442 49698
rect 31442 49646 31444 49698
rect 31388 49644 31444 49646
rect 29260 49532 29316 49588
rect 27468 48748 27524 48804
rect 27916 47682 27972 47684
rect 27916 47630 27918 47682
rect 27918 47630 27970 47682
rect 27970 47630 27972 47682
rect 27916 47628 27972 47630
rect 26908 47292 26964 47348
rect 26908 46844 26964 46900
rect 34412 49810 34468 49812
rect 34412 49758 34414 49810
rect 34414 49758 34466 49810
rect 34466 49758 34468 49810
rect 34412 49756 34468 49758
rect 34748 49756 34804 49812
rect 33964 48748 34020 48804
rect 33404 48076 33460 48132
rect 31948 47292 32004 47348
rect 28252 47180 28308 47236
rect 31164 47234 31220 47236
rect 31164 47182 31166 47234
rect 31166 47182 31218 47234
rect 31218 47182 31220 47234
rect 31164 47180 31220 47182
rect 28028 46732 28084 46788
rect 30044 46786 30100 46788
rect 30044 46734 30046 46786
rect 30046 46734 30098 46786
rect 30098 46734 30100 46786
rect 30044 46732 30100 46734
rect 26348 45666 26404 45668
rect 26348 45614 26350 45666
rect 26350 45614 26402 45666
rect 26402 45614 26404 45666
rect 26348 45612 26404 45614
rect 26124 43596 26180 43652
rect 26572 43596 26628 43652
rect 25004 42754 25060 42756
rect 25004 42702 25006 42754
rect 25006 42702 25058 42754
rect 25058 42702 25060 42754
rect 25004 42700 25060 42702
rect 25340 42700 25396 42756
rect 23884 42588 23940 42644
rect 21980 42252 22036 42308
rect 22428 42252 22484 42308
rect 24444 42642 24500 42644
rect 24444 42590 24446 42642
rect 24446 42590 24498 42642
rect 24498 42590 24500 42642
rect 24444 42588 24500 42590
rect 25228 42642 25284 42644
rect 25228 42590 25230 42642
rect 25230 42590 25282 42642
rect 25282 42590 25284 42642
rect 25228 42588 25284 42590
rect 23212 41970 23268 41972
rect 23212 41918 23214 41970
rect 23214 41918 23266 41970
rect 23266 41918 23268 41970
rect 23212 41916 23268 41918
rect 23100 41692 23156 41748
rect 24556 41970 24612 41972
rect 24556 41918 24558 41970
rect 24558 41918 24610 41970
rect 24610 41918 24612 41970
rect 24556 41916 24612 41918
rect 24220 41804 24276 41860
rect 23996 41692 24052 41748
rect 22652 41186 22708 41188
rect 22652 41134 22654 41186
rect 22654 41134 22706 41186
rect 22706 41134 22708 41186
rect 22652 41132 22708 41134
rect 22428 40348 22484 40404
rect 21644 39730 21700 39732
rect 21644 39678 21646 39730
rect 21646 39678 21698 39730
rect 21698 39678 21700 39730
rect 21644 39676 21700 39678
rect 22092 39676 22148 39732
rect 20972 39228 21028 39284
rect 22092 39228 22148 39284
rect 26348 42866 26404 42868
rect 26348 42814 26350 42866
rect 26350 42814 26402 42866
rect 26402 42814 26404 42866
rect 26348 42812 26404 42814
rect 26684 42866 26740 42868
rect 26684 42814 26686 42866
rect 26686 42814 26738 42866
rect 26738 42814 26740 42866
rect 26684 42812 26740 42814
rect 25788 42194 25844 42196
rect 25788 42142 25790 42194
rect 25790 42142 25842 42194
rect 25842 42142 25844 42194
rect 25788 42140 25844 42142
rect 25116 41970 25172 41972
rect 25116 41918 25118 41970
rect 25118 41918 25170 41970
rect 25170 41918 25172 41970
rect 25116 41916 25172 41918
rect 25340 39394 25396 39396
rect 25340 39342 25342 39394
rect 25342 39342 25394 39394
rect 25394 39342 25396 39394
rect 25340 39340 25396 39342
rect 25452 39004 25508 39060
rect 20412 35698 20468 35700
rect 20412 35646 20414 35698
rect 20414 35646 20466 35698
rect 20466 35646 20468 35698
rect 20412 35644 20468 35646
rect 20524 34972 20580 35028
rect 19180 31612 19236 31668
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20412 31106 20468 31108
rect 20412 31054 20414 31106
rect 20414 31054 20466 31106
rect 20466 31054 20468 31106
rect 20412 31052 20468 31054
rect 18284 30882 18340 30884
rect 18284 30830 18286 30882
rect 18286 30830 18338 30882
rect 18338 30830 18340 30882
rect 18284 30828 18340 30830
rect 17948 30322 18004 30324
rect 17948 30270 17950 30322
rect 17950 30270 18002 30322
rect 18002 30270 18004 30322
rect 17948 30268 18004 30270
rect 18172 30210 18228 30212
rect 18172 30158 18174 30210
rect 18174 30158 18226 30210
rect 18226 30158 18228 30210
rect 18172 30156 18228 30158
rect 19404 30268 19460 30324
rect 17724 29260 17780 29316
rect 17724 29036 17780 29092
rect 17612 28642 17668 28644
rect 17612 28590 17614 28642
rect 17614 28590 17666 28642
rect 17666 28590 17668 28642
rect 17612 28588 17668 28590
rect 16828 24780 16884 24836
rect 16716 24668 16772 24724
rect 15932 22594 15988 22596
rect 15932 22542 15934 22594
rect 15934 22542 15986 22594
rect 15986 22542 15988 22594
rect 15932 22540 15988 22542
rect 16716 20636 16772 20692
rect 16828 21532 16884 21588
rect 18844 29260 18900 29316
rect 18172 28700 18228 28756
rect 18732 28754 18788 28756
rect 18732 28702 18734 28754
rect 18734 28702 18786 28754
rect 18786 28702 18788 28754
rect 18732 28700 18788 28702
rect 19068 27858 19124 27860
rect 19068 27806 19070 27858
rect 19070 27806 19122 27858
rect 19122 27806 19124 27858
rect 19068 27804 19124 27806
rect 18284 26124 18340 26180
rect 18396 25676 18452 25732
rect 17948 25506 18004 25508
rect 17948 25454 17950 25506
rect 17950 25454 18002 25506
rect 18002 25454 18004 25506
rect 17948 25452 18004 25454
rect 18396 25228 18452 25284
rect 18844 26178 18900 26180
rect 18844 26126 18846 26178
rect 18846 26126 18898 26178
rect 18898 26126 18900 26178
rect 18844 26124 18900 26126
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 28924 19684 28980
rect 20076 28700 20132 28756
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 28028 19684 28084
rect 20300 28028 20356 28084
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 25730 19684 25732
rect 19628 25678 19630 25730
rect 19630 25678 19682 25730
rect 19682 25678 19684 25730
rect 19628 25676 19684 25678
rect 18620 25506 18676 25508
rect 18620 25454 18622 25506
rect 18622 25454 18674 25506
rect 18674 25454 18676 25506
rect 18620 25452 18676 25454
rect 19068 25228 19124 25284
rect 18956 24892 19012 24948
rect 18284 24722 18340 24724
rect 18284 24670 18286 24722
rect 18286 24670 18338 24722
rect 18338 24670 18340 24722
rect 18284 24668 18340 24670
rect 19068 24780 19124 24836
rect 19516 25506 19572 25508
rect 19516 25454 19518 25506
rect 19518 25454 19570 25506
rect 19570 25454 19572 25506
rect 19516 25452 19572 25454
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24892 20244 24948
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18508 23324 18564 23380
rect 18284 23212 18340 23268
rect 19516 23154 19572 23156
rect 19516 23102 19518 23154
rect 19518 23102 19570 23154
rect 19570 23102 19572 23154
rect 19516 23100 19572 23102
rect 21980 35196 22036 35252
rect 21980 33964 22036 34020
rect 22428 34188 22484 34244
rect 21980 32562 22036 32564
rect 21980 32510 21982 32562
rect 21982 32510 22034 32562
rect 22034 32510 22036 32562
rect 21980 32508 22036 32510
rect 21868 31724 21924 31780
rect 21532 31612 21588 31668
rect 21084 31164 21140 31220
rect 20748 28754 20804 28756
rect 20748 28702 20750 28754
rect 20750 28702 20802 28754
rect 20802 28702 20804 28754
rect 20748 28700 20804 28702
rect 20972 28140 21028 28196
rect 21084 29820 21140 29876
rect 20636 28028 20692 28084
rect 20636 26572 20692 26628
rect 20524 23212 20580 23268
rect 20412 23100 20468 23156
rect 18956 22258 19012 22260
rect 18956 22206 18958 22258
rect 18958 22206 19010 22258
rect 19010 22206 19012 22258
rect 18956 22204 19012 22206
rect 20636 22204 20692 22260
rect 17724 22146 17780 22148
rect 17724 22094 17726 22146
rect 17726 22094 17778 22146
rect 17778 22094 17780 22146
rect 17724 22092 17780 22094
rect 18620 22146 18676 22148
rect 18620 22094 18622 22146
rect 18622 22094 18674 22146
rect 18674 22094 18676 22146
rect 18620 22092 18676 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 17724 21586 17780 21588
rect 17724 21534 17726 21586
rect 17726 21534 17778 21586
rect 17778 21534 17780 21586
rect 17724 21532 17780 21534
rect 17500 21308 17556 21364
rect 18284 21308 18340 21364
rect 16604 20578 16660 20580
rect 16604 20526 16606 20578
rect 16606 20526 16658 20578
rect 16658 20526 16660 20578
rect 16604 20524 16660 20526
rect 16044 20412 16100 20468
rect 15708 20130 15764 20132
rect 15708 20078 15710 20130
rect 15710 20078 15762 20130
rect 15762 20078 15764 20130
rect 15708 20076 15764 20078
rect 15484 19964 15540 20020
rect 16044 19852 16100 19908
rect 16268 19906 16324 19908
rect 16268 19854 16270 19906
rect 16270 19854 16322 19906
rect 16322 19854 16324 19906
rect 16268 19852 16324 19854
rect 15372 18508 15428 18564
rect 16268 18450 16324 18452
rect 16268 18398 16270 18450
rect 16270 18398 16322 18450
rect 16322 18398 16324 18450
rect 16268 18396 16324 18398
rect 15932 18284 15988 18340
rect 15484 17164 15540 17220
rect 15820 17106 15876 17108
rect 15820 17054 15822 17106
rect 15822 17054 15874 17106
rect 15874 17054 15876 17106
rect 15820 17052 15876 17054
rect 16380 17388 16436 17444
rect 15820 15932 15876 15988
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 17500 19852 17556 19908
rect 17052 19346 17108 19348
rect 17052 19294 17054 19346
rect 17054 19294 17106 19346
rect 17106 19294 17108 19346
rect 17052 19292 17108 19294
rect 17052 17442 17108 17444
rect 17052 17390 17054 17442
rect 17054 17390 17106 17442
rect 17106 17390 17108 17442
rect 17052 17388 17108 17390
rect 20300 19628 20356 19684
rect 20524 19740 20580 19796
rect 18172 19292 18228 19348
rect 20412 19404 20468 19460
rect 20188 19010 20244 19012
rect 20188 18958 20190 19010
rect 20190 18958 20242 19010
rect 20242 18958 20244 19010
rect 20188 18956 20244 18958
rect 16492 17052 16548 17108
rect 17612 17164 17668 17220
rect 16156 16770 16212 16772
rect 16156 16718 16158 16770
rect 16158 16718 16210 16770
rect 16210 16718 16212 16770
rect 16156 16716 16212 16718
rect 16492 16658 16548 16660
rect 16492 16606 16494 16658
rect 16494 16606 16546 16658
rect 16546 16606 16548 16658
rect 16492 16604 16548 16606
rect 16604 16268 16660 16324
rect 17948 17052 18004 17108
rect 16716 16044 16772 16100
rect 17276 16828 17332 16884
rect 17500 16828 17556 16884
rect 15148 14530 15204 14532
rect 15148 14478 15150 14530
rect 15150 14478 15202 14530
rect 15202 14478 15204 14530
rect 15148 14476 15204 14478
rect 14364 13804 14420 13860
rect 13916 13132 13972 13188
rect 13468 12738 13524 12740
rect 13468 12686 13470 12738
rect 13470 12686 13522 12738
rect 13522 12686 13524 12738
rect 13468 12684 13524 12686
rect 10668 11282 10724 11284
rect 10668 11230 10670 11282
rect 10670 11230 10722 11282
rect 10722 11230 10724 11282
rect 10668 11228 10724 11230
rect 9660 8876 9716 8932
rect 10668 10610 10724 10612
rect 10668 10558 10670 10610
rect 10670 10558 10722 10610
rect 10722 10558 10724 10610
rect 10668 10556 10724 10558
rect 11116 11618 11172 11620
rect 11116 11566 11118 11618
rect 11118 11566 11170 11618
rect 11170 11566 11172 11618
rect 11116 11564 11172 11566
rect 12796 11394 12852 11396
rect 12796 11342 12798 11394
rect 12798 11342 12850 11394
rect 12850 11342 12852 11394
rect 12796 11340 12852 11342
rect 13468 11394 13524 11396
rect 13468 11342 13470 11394
rect 13470 11342 13522 11394
rect 13522 11342 13524 11394
rect 13468 11340 13524 11342
rect 11116 10610 11172 10612
rect 11116 10558 11118 10610
rect 11118 10558 11170 10610
rect 11170 10558 11172 10610
rect 11116 10556 11172 10558
rect 11116 9996 11172 10052
rect 11564 9884 11620 9940
rect 12460 10444 12516 10500
rect 12348 9996 12404 10052
rect 12908 10668 12964 10724
rect 13468 10444 13524 10500
rect 14140 13356 14196 13412
rect 14588 13356 14644 13412
rect 14028 11564 14084 11620
rect 13916 10722 13972 10724
rect 13916 10670 13918 10722
rect 13918 10670 13970 10722
rect 13970 10670 13972 10722
rect 13916 10668 13972 10670
rect 15148 12684 15204 12740
rect 16044 15932 16100 15988
rect 15708 14530 15764 14532
rect 15708 14478 15710 14530
rect 15710 14478 15762 14530
rect 15762 14478 15764 14530
rect 15708 14476 15764 14478
rect 15372 14418 15428 14420
rect 15372 14366 15374 14418
rect 15374 14366 15426 14418
rect 15426 14366 15428 14418
rect 15372 14364 15428 14366
rect 17388 16268 17444 16324
rect 17276 15986 17332 15988
rect 17276 15934 17278 15986
rect 17278 15934 17330 15986
rect 17330 15934 17332 15986
rect 17276 15932 17332 15934
rect 17836 16770 17892 16772
rect 17836 16718 17838 16770
rect 17838 16718 17890 16770
rect 17890 16718 17892 16770
rect 17836 16716 17892 16718
rect 19068 16716 19124 16772
rect 18172 15538 18228 15540
rect 18172 15486 18174 15538
rect 18174 15486 18226 15538
rect 18226 15486 18228 15538
rect 18172 15484 18228 15486
rect 17388 14530 17444 14532
rect 17388 14478 17390 14530
rect 17390 14478 17442 14530
rect 17442 14478 17444 14530
rect 17388 14476 17444 14478
rect 16044 14306 16100 14308
rect 16044 14254 16046 14306
rect 16046 14254 16098 14306
rect 16098 14254 16100 14306
rect 16044 14252 16100 14254
rect 16380 14364 16436 14420
rect 15932 13186 15988 13188
rect 15932 13134 15934 13186
rect 15934 13134 15986 13186
rect 15986 13134 15988 13186
rect 15932 13132 15988 13134
rect 15260 12572 15316 12628
rect 15148 12012 15204 12068
rect 14924 10668 14980 10724
rect 15036 11564 15092 11620
rect 12684 9884 12740 9940
rect 11788 9826 11844 9828
rect 11788 9774 11790 9826
rect 11790 9774 11842 9826
rect 11842 9774 11844 9826
rect 11788 9772 11844 9774
rect 11004 9602 11060 9604
rect 11004 9550 11006 9602
rect 11006 9550 11058 9602
rect 11058 9550 11060 9602
rect 11004 9548 11060 9550
rect 11228 9548 11284 9604
rect 12124 9602 12180 9604
rect 12124 9550 12126 9602
rect 12126 9550 12178 9602
rect 12178 9550 12180 9602
rect 12124 9548 12180 9550
rect 12684 9714 12740 9716
rect 12684 9662 12686 9714
rect 12686 9662 12738 9714
rect 12738 9662 12740 9714
rect 12684 9660 12740 9662
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 8988 6636 9044 6692
rect 9100 6466 9156 6468
rect 9100 6414 9102 6466
rect 9102 6414 9154 6466
rect 9154 6414 9156 6466
rect 9100 6412 9156 6414
rect 13244 9884 13300 9940
rect 12908 9826 12964 9828
rect 12908 9774 12910 9826
rect 12910 9774 12962 9826
rect 12962 9774 12964 9826
rect 12908 9772 12964 9774
rect 13916 9884 13972 9940
rect 17164 14418 17220 14420
rect 17164 14366 17166 14418
rect 17166 14366 17218 14418
rect 17218 14366 17220 14418
rect 17164 14364 17220 14366
rect 17388 13020 17444 13076
rect 16156 12850 16212 12852
rect 16156 12798 16158 12850
rect 16158 12798 16210 12850
rect 16210 12798 16212 12850
rect 16156 12796 16212 12798
rect 16828 12850 16884 12852
rect 16828 12798 16830 12850
rect 16830 12798 16882 12850
rect 16882 12798 16884 12850
rect 16828 12796 16884 12798
rect 15820 12178 15876 12180
rect 15820 12126 15822 12178
rect 15822 12126 15874 12178
rect 15874 12126 15876 12178
rect 15820 12124 15876 12126
rect 16044 12684 16100 12740
rect 15260 10556 15316 10612
rect 15148 9884 15204 9940
rect 14476 9826 14532 9828
rect 14476 9774 14478 9826
rect 14478 9774 14530 9826
rect 14530 9774 14532 9826
rect 14476 9772 14532 9774
rect 13580 9660 13636 9716
rect 14252 9548 14308 9604
rect 14700 9660 14756 9716
rect 10220 7474 10276 7476
rect 10220 7422 10222 7474
rect 10222 7422 10274 7474
rect 10274 7422 10276 7474
rect 10220 7420 10276 7422
rect 10668 7420 10724 7476
rect 13580 7362 13636 7364
rect 13580 7310 13582 7362
rect 13582 7310 13634 7362
rect 13634 7310 13636 7362
rect 13580 7308 13636 7310
rect 9884 6636 9940 6692
rect 10668 6748 10724 6804
rect 12348 6636 12404 6692
rect 10556 6466 10612 6468
rect 10556 6414 10558 6466
rect 10558 6414 10610 6466
rect 10610 6414 10612 6466
rect 10556 6412 10612 6414
rect 10556 5180 10612 5236
rect 11900 5234 11956 5236
rect 11900 5182 11902 5234
rect 11902 5182 11954 5234
rect 11954 5182 11956 5234
rect 11900 5180 11956 5182
rect 13468 6690 13524 6692
rect 13468 6638 13470 6690
rect 13470 6638 13522 6690
rect 13522 6638 13524 6690
rect 13468 6636 13524 6638
rect 14588 7308 14644 7364
rect 15820 11116 15876 11172
rect 15372 9772 15428 9828
rect 16380 12236 16436 12292
rect 17724 14364 17780 14420
rect 18844 15314 18900 15316
rect 18844 15262 18846 15314
rect 18846 15262 18898 15314
rect 18898 15262 18900 15314
rect 18844 15260 18900 15262
rect 17612 13186 17668 13188
rect 17612 13134 17614 13186
rect 17614 13134 17666 13186
rect 17666 13134 17668 13186
rect 17612 13132 17668 13134
rect 17948 13468 18004 13524
rect 17836 12962 17892 12964
rect 17836 12910 17838 12962
rect 17838 12910 17890 12962
rect 17890 12910 17892 12962
rect 17836 12908 17892 12910
rect 16828 10610 16884 10612
rect 16828 10558 16830 10610
rect 16830 10558 16882 10610
rect 16882 10558 16884 10610
rect 16828 10556 16884 10558
rect 19516 15484 19572 15540
rect 19068 14530 19124 14532
rect 19068 14478 19070 14530
rect 19070 14478 19122 14530
rect 19122 14478 19124 14530
rect 19068 14476 19124 14478
rect 18396 14418 18452 14420
rect 18396 14366 18398 14418
rect 18398 14366 18450 14418
rect 18450 14366 18452 14418
rect 18396 14364 18452 14366
rect 18284 14252 18340 14308
rect 18508 13468 18564 13524
rect 19068 13132 19124 13188
rect 18396 12962 18452 12964
rect 18396 12910 18398 12962
rect 18398 12910 18450 12962
rect 18450 12910 18452 12962
rect 18396 12908 18452 12910
rect 18060 12236 18116 12292
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 16882 20132 16884
rect 20076 16830 20078 16882
rect 20078 16830 20130 16882
rect 20130 16830 20132 16882
rect 20076 16828 20132 16830
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20300 15036 20356 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 18620 12124 18676 12180
rect 17724 11676 17780 11732
rect 17500 10556 17556 10612
rect 20300 11564 20356 11620
rect 21644 31106 21700 31108
rect 21644 31054 21646 31106
rect 21646 31054 21698 31106
rect 21698 31054 21700 31106
rect 21644 31052 21700 31054
rect 21532 30994 21588 30996
rect 21532 30942 21534 30994
rect 21534 30942 21586 30994
rect 21586 30942 21588 30994
rect 21532 30940 21588 30942
rect 22876 36428 22932 36484
rect 22652 36370 22708 36372
rect 22652 36318 22654 36370
rect 22654 36318 22706 36370
rect 22706 36318 22708 36370
rect 22652 36316 22708 36318
rect 25340 36482 25396 36484
rect 25340 36430 25342 36482
rect 25342 36430 25394 36482
rect 25394 36430 25396 36482
rect 25340 36428 25396 36430
rect 24332 36370 24388 36372
rect 24332 36318 24334 36370
rect 24334 36318 24386 36370
rect 24386 36318 24388 36370
rect 24332 36316 24388 36318
rect 23100 35420 23156 35476
rect 23436 35196 23492 35252
rect 24220 35420 24276 35476
rect 25340 35308 25396 35364
rect 24220 34972 24276 35028
rect 25676 37436 25732 37492
rect 26124 42028 26180 42084
rect 26348 41970 26404 41972
rect 26348 41918 26350 41970
rect 26350 41918 26402 41970
rect 26402 41918 26404 41970
rect 26348 41916 26404 41918
rect 26124 37378 26180 37380
rect 26124 37326 26126 37378
rect 26126 37326 26178 37378
rect 26178 37326 26180 37378
rect 26124 37324 26180 37326
rect 25788 35698 25844 35700
rect 25788 35646 25790 35698
rect 25790 35646 25842 35698
rect 25842 35646 25844 35698
rect 25788 35644 25844 35646
rect 26796 35698 26852 35700
rect 26796 35646 26798 35698
rect 26798 35646 26850 35698
rect 26850 35646 26852 35698
rect 26796 35644 26852 35646
rect 27804 45836 27860 45892
rect 27020 42812 27076 42868
rect 27468 42530 27524 42532
rect 27468 42478 27470 42530
rect 27470 42478 27522 42530
rect 27522 42478 27524 42530
rect 27468 42476 27524 42478
rect 27468 42028 27524 42084
rect 28812 45218 28868 45220
rect 28812 45166 28814 45218
rect 28814 45166 28866 45218
rect 28866 45166 28868 45218
rect 28812 45164 28868 45166
rect 28140 44940 28196 44996
rect 27916 42754 27972 42756
rect 27916 42702 27918 42754
rect 27918 42702 27970 42754
rect 27970 42702 27972 42754
rect 27916 42700 27972 42702
rect 27692 39564 27748 39620
rect 29260 45052 29316 45108
rect 28364 43596 28420 43652
rect 28364 42924 28420 42980
rect 28364 39618 28420 39620
rect 28364 39566 28366 39618
rect 28366 39566 28418 39618
rect 28418 39566 28420 39618
rect 28364 39564 28420 39566
rect 29596 45106 29652 45108
rect 29596 45054 29598 45106
rect 29598 45054 29650 45106
rect 29650 45054 29652 45106
rect 29596 45052 29652 45054
rect 30716 45052 30772 45108
rect 28812 43650 28868 43652
rect 28812 43598 28814 43650
rect 28814 43598 28866 43650
rect 28866 43598 28868 43650
rect 28812 43596 28868 43598
rect 29260 42754 29316 42756
rect 29260 42702 29262 42754
rect 29262 42702 29314 42754
rect 29314 42702 29316 42754
rect 29260 42700 29316 42702
rect 28588 42530 28644 42532
rect 28588 42478 28590 42530
rect 28590 42478 28642 42530
rect 28642 42478 28644 42530
rect 28588 42476 28644 42478
rect 29708 42754 29764 42756
rect 29708 42702 29710 42754
rect 29710 42702 29762 42754
rect 29762 42702 29764 42754
rect 29708 42700 29764 42702
rect 29484 42476 29540 42532
rect 31500 43260 31556 43316
rect 31388 42924 31444 42980
rect 29820 41970 29876 41972
rect 29820 41918 29822 41970
rect 29822 41918 29874 41970
rect 29874 41918 29876 41970
rect 29820 41916 29876 41918
rect 29148 41858 29204 41860
rect 29148 41806 29150 41858
rect 29150 41806 29202 41858
rect 29202 41806 29204 41858
rect 29148 41804 29204 41806
rect 27020 38556 27076 38612
rect 27020 37772 27076 37828
rect 27916 38332 27972 38388
rect 28476 38556 28532 38612
rect 28588 38220 28644 38276
rect 28588 38050 28644 38052
rect 28588 37998 28590 38050
rect 28590 37998 28642 38050
rect 28642 37998 28644 38050
rect 28588 37996 28644 37998
rect 27132 35868 27188 35924
rect 24668 34748 24724 34804
rect 24332 34242 24388 34244
rect 24332 34190 24334 34242
rect 24334 34190 24386 34242
rect 24386 34190 24388 34242
rect 24332 34188 24388 34190
rect 22652 32508 22708 32564
rect 22204 31052 22260 31108
rect 22316 30994 22372 30996
rect 22316 30942 22318 30994
rect 22318 30942 22370 30994
rect 22370 30942 22372 30994
rect 22316 30940 22372 30942
rect 22764 31164 22820 31220
rect 22540 30828 22596 30884
rect 21756 30156 21812 30212
rect 22316 30210 22372 30212
rect 22316 30158 22318 30210
rect 22318 30158 22370 30210
rect 22370 30158 22372 30210
rect 22316 30156 22372 30158
rect 21980 29820 22036 29876
rect 21868 28476 21924 28532
rect 22540 30098 22596 30100
rect 22540 30046 22542 30098
rect 22542 30046 22594 30098
rect 22594 30046 22596 30098
rect 22540 30044 22596 30046
rect 22652 29596 22708 29652
rect 22652 28700 22708 28756
rect 22540 28530 22596 28532
rect 22540 28478 22542 28530
rect 22542 28478 22594 28530
rect 22594 28478 22596 28530
rect 22540 28476 22596 28478
rect 22428 27804 22484 27860
rect 21980 27580 22036 27636
rect 22652 28028 22708 28084
rect 24892 33458 24948 33460
rect 24892 33406 24894 33458
rect 24894 33406 24946 33458
rect 24946 33406 24948 33458
rect 24892 33404 24948 33406
rect 24780 33292 24836 33348
rect 24332 32844 24388 32900
rect 23548 31724 23604 31780
rect 22988 31052 23044 31108
rect 23100 30098 23156 30100
rect 23100 30046 23102 30098
rect 23102 30046 23154 30098
rect 23154 30046 23156 30098
rect 23100 30044 23156 30046
rect 22876 29260 22932 29316
rect 23212 28754 23268 28756
rect 23212 28702 23214 28754
rect 23214 28702 23266 28754
rect 23266 28702 23268 28754
rect 23212 28700 23268 28702
rect 22316 27020 22372 27076
rect 21644 26908 21700 26964
rect 22204 26962 22260 26964
rect 22204 26910 22206 26962
rect 22206 26910 22258 26962
rect 22258 26910 22260 26962
rect 22204 26908 22260 26910
rect 22540 26962 22596 26964
rect 22540 26910 22542 26962
rect 22542 26910 22594 26962
rect 22594 26910 22596 26962
rect 22540 26908 22596 26910
rect 23212 28364 23268 28420
rect 23660 31612 23716 31668
rect 23884 30828 23940 30884
rect 24108 30156 24164 30212
rect 23772 29484 23828 29540
rect 23324 27580 23380 27636
rect 23212 27132 23268 27188
rect 23884 27186 23940 27188
rect 23884 27134 23886 27186
rect 23886 27134 23938 27186
rect 23938 27134 23940 27186
rect 23884 27132 23940 27134
rect 21644 25676 21700 25732
rect 22316 25676 22372 25732
rect 21308 24892 21364 24948
rect 22540 24780 22596 24836
rect 21196 23154 21252 23156
rect 21196 23102 21198 23154
rect 21198 23102 21250 23154
rect 21250 23102 21252 23154
rect 21196 23100 21252 23102
rect 21308 21474 21364 21476
rect 21308 21422 21310 21474
rect 21310 21422 21362 21474
rect 21362 21422 21364 21474
rect 21308 21420 21364 21422
rect 21420 19906 21476 19908
rect 21420 19854 21422 19906
rect 21422 19854 21474 19906
rect 21474 19854 21476 19906
rect 21420 19852 21476 19854
rect 22988 24722 23044 24724
rect 22988 24670 22990 24722
rect 22990 24670 23042 24722
rect 23042 24670 23044 24722
rect 22988 24668 23044 24670
rect 23660 24668 23716 24724
rect 23660 22316 23716 22372
rect 24108 27970 24164 27972
rect 24108 27918 24110 27970
rect 24110 27918 24162 27970
rect 24162 27918 24164 27970
rect 24108 27916 24164 27918
rect 24220 27858 24276 27860
rect 24220 27806 24222 27858
rect 24222 27806 24274 27858
rect 24274 27806 24276 27858
rect 24220 27804 24276 27806
rect 25004 31612 25060 31668
rect 25004 30210 25060 30212
rect 25004 30158 25006 30210
rect 25006 30158 25058 30210
rect 25058 30158 25060 30210
rect 25004 30156 25060 30158
rect 24444 26290 24500 26292
rect 24444 26238 24446 26290
rect 24446 26238 24498 26290
rect 24498 26238 24500 26290
rect 24444 26236 24500 26238
rect 23996 21586 24052 21588
rect 23996 21534 23998 21586
rect 23998 21534 24050 21586
rect 24050 21534 24052 21586
rect 23996 21532 24052 21534
rect 23548 21420 23604 21476
rect 22764 17388 22820 17444
rect 24332 22370 24388 22372
rect 24332 22318 24334 22370
rect 24334 22318 24386 22370
rect 24386 22318 24388 22370
rect 24332 22316 24388 22318
rect 24220 21532 24276 21588
rect 24668 28252 24724 28308
rect 24668 27916 24724 27972
rect 24780 24050 24836 24052
rect 24780 23998 24782 24050
rect 24782 23998 24834 24050
rect 24834 23998 24836 24050
rect 24780 23996 24836 23998
rect 24556 21644 24612 21700
rect 24780 23100 24836 23156
rect 24108 20300 24164 20356
rect 23100 19404 23156 19460
rect 21084 16716 21140 16772
rect 21644 16770 21700 16772
rect 21644 16718 21646 16770
rect 21646 16718 21698 16770
rect 21698 16718 21700 16770
rect 21644 16716 21700 16718
rect 23324 18956 23380 19012
rect 23436 17948 23492 18004
rect 23100 16098 23156 16100
rect 23100 16046 23102 16098
rect 23102 16046 23154 16098
rect 23154 16046 23156 16098
rect 23100 16044 23156 16046
rect 23324 16716 23380 16772
rect 20972 15260 21028 15316
rect 22092 15314 22148 15316
rect 22092 15262 22094 15314
rect 22094 15262 22146 15314
rect 22146 15262 22148 15314
rect 22092 15260 22148 15262
rect 21756 13634 21812 13636
rect 21756 13582 21758 13634
rect 21758 13582 21810 13634
rect 21810 13582 21812 13634
rect 21756 13580 21812 13582
rect 20860 13522 20916 13524
rect 20860 13470 20862 13522
rect 20862 13470 20914 13522
rect 20914 13470 20916 13522
rect 20860 13468 20916 13470
rect 22876 12684 22932 12740
rect 19628 11116 19684 11172
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 16156 9772 16212 9828
rect 16716 9548 16772 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 9100 19684 9156
rect 23884 19852 23940 19908
rect 24780 19964 24836 20020
rect 24108 19292 24164 19348
rect 24444 19292 24500 19348
rect 23996 19234 24052 19236
rect 23996 19182 23998 19234
rect 23998 19182 24050 19234
rect 24050 19182 24052 19234
rect 23996 19180 24052 19182
rect 24332 18956 24388 19012
rect 24332 17500 24388 17556
rect 23772 17052 23828 17108
rect 24220 17106 24276 17108
rect 24220 17054 24222 17106
rect 24222 17054 24274 17106
rect 24274 17054 24276 17106
rect 24220 17052 24276 17054
rect 24108 16716 24164 16772
rect 24556 19180 24612 19236
rect 25004 22258 25060 22260
rect 25004 22206 25006 22258
rect 25006 22206 25058 22258
rect 25058 22206 25060 22258
rect 25004 22204 25060 22206
rect 25676 34802 25732 34804
rect 25676 34750 25678 34802
rect 25678 34750 25730 34802
rect 25730 34750 25732 34802
rect 25676 34748 25732 34750
rect 27132 35308 27188 35364
rect 25564 33404 25620 33460
rect 25452 32562 25508 32564
rect 25452 32510 25454 32562
rect 25454 32510 25506 32562
rect 25506 32510 25508 32562
rect 25452 32508 25508 32510
rect 26236 33180 26292 33236
rect 25564 32396 25620 32452
rect 26012 31554 26068 31556
rect 26012 31502 26014 31554
rect 26014 31502 26066 31554
rect 26066 31502 26068 31554
rect 26012 31500 26068 31502
rect 25452 31052 25508 31108
rect 26012 30268 26068 30324
rect 26348 32508 26404 32564
rect 27132 33964 27188 34020
rect 27020 33234 27076 33236
rect 27020 33182 27022 33234
rect 27022 33182 27074 33234
rect 27074 33182 27076 33234
rect 27020 33180 27076 33182
rect 26460 31554 26516 31556
rect 26460 31502 26462 31554
rect 26462 31502 26514 31554
rect 26514 31502 26516 31554
rect 26460 31500 26516 31502
rect 26684 31276 26740 31332
rect 28252 33964 28308 34020
rect 29372 41804 29428 41860
rect 29260 39564 29316 39620
rect 30380 41916 30436 41972
rect 31052 41074 31108 41076
rect 31052 41022 31054 41074
rect 31054 41022 31106 41074
rect 31106 41022 31108 41074
rect 31052 41020 31108 41022
rect 30044 40626 30100 40628
rect 30044 40574 30046 40626
rect 30046 40574 30098 40626
rect 30098 40574 30100 40626
rect 30044 40572 30100 40574
rect 30716 40626 30772 40628
rect 30716 40574 30718 40626
rect 30718 40574 30770 40626
rect 30770 40574 30772 40626
rect 30716 40572 30772 40574
rect 33180 47180 33236 47236
rect 31724 42924 31780 42980
rect 31948 44380 32004 44436
rect 32060 44492 32116 44548
rect 33068 45218 33124 45220
rect 33068 45166 33070 45218
rect 33070 45166 33122 45218
rect 33122 45166 33124 45218
rect 33068 45164 33124 45166
rect 32396 45106 32452 45108
rect 32396 45054 32398 45106
rect 32398 45054 32450 45106
rect 32450 45054 32452 45106
rect 32396 45052 32452 45054
rect 33516 44828 33572 44884
rect 33852 45052 33908 45108
rect 33852 44492 33908 44548
rect 32732 44380 32788 44436
rect 32396 44322 32452 44324
rect 32396 44270 32398 44322
rect 32398 44270 32450 44322
rect 32450 44270 32452 44322
rect 32396 44268 32452 44270
rect 32172 43372 32228 43428
rect 32060 43314 32116 43316
rect 32060 43262 32062 43314
rect 32062 43262 32114 43314
rect 32114 43262 32116 43314
rect 32060 43260 32116 43262
rect 32396 43260 32452 43316
rect 32060 42812 32116 42868
rect 33628 44322 33684 44324
rect 33628 44270 33630 44322
rect 33630 44270 33682 44322
rect 33682 44270 33684 44322
rect 33628 44268 33684 44270
rect 33516 44156 33572 44212
rect 32732 42866 32788 42868
rect 32732 42814 32734 42866
rect 32734 42814 32786 42866
rect 32786 42814 32788 42866
rect 32732 42812 32788 42814
rect 36764 50034 36820 50036
rect 36764 49982 36766 50034
rect 36766 49982 36818 50034
rect 36818 49982 36820 50034
rect 36764 49980 36820 49982
rect 37212 49980 37268 50036
rect 39116 50482 39172 50484
rect 39116 50430 39118 50482
rect 39118 50430 39170 50482
rect 39170 50430 39172 50482
rect 39116 50428 39172 50430
rect 39788 49980 39844 50036
rect 41020 50428 41076 50484
rect 37772 49922 37828 49924
rect 37772 49870 37774 49922
rect 37774 49870 37826 49922
rect 37826 49870 37828 49922
rect 37772 49868 37828 49870
rect 36652 49810 36708 49812
rect 36652 49758 36654 49810
rect 36654 49758 36706 49810
rect 36706 49758 36708 49810
rect 36652 49756 36708 49758
rect 36876 49698 36932 49700
rect 36876 49646 36878 49698
rect 36878 49646 36930 49698
rect 36930 49646 36932 49698
rect 36876 49644 36932 49646
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 48748 35140 48804
rect 34860 48636 34916 48692
rect 39004 49756 39060 49812
rect 37548 49698 37604 49700
rect 37548 49646 37550 49698
rect 37550 49646 37602 49698
rect 37602 49646 37604 49698
rect 37548 49644 37604 49646
rect 37772 48860 37828 48916
rect 36988 48636 37044 48692
rect 34300 48188 34356 48244
rect 34188 44492 34244 44548
rect 34188 43820 34244 43876
rect 34188 43148 34244 43204
rect 33628 42476 33684 42532
rect 31948 41804 32004 41860
rect 34524 48130 34580 48132
rect 34524 48078 34526 48130
rect 34526 48078 34578 48130
rect 34578 48078 34580 48130
rect 34524 48076 34580 48078
rect 34972 48242 35028 48244
rect 34972 48190 34974 48242
rect 34974 48190 35026 48242
rect 35026 48190 35028 48242
rect 34972 48188 35028 48190
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 47346 35252 47348
rect 35196 47294 35198 47346
rect 35198 47294 35250 47346
rect 35250 47294 35252 47346
rect 35196 47292 35252 47294
rect 37772 47682 37828 47684
rect 37772 47630 37774 47682
rect 37774 47630 37826 47682
rect 37826 47630 37828 47682
rect 37772 47628 37828 47630
rect 34412 43596 34468 43652
rect 34860 44994 34916 44996
rect 34860 44942 34862 44994
rect 34862 44942 34914 44994
rect 34914 44942 34916 44994
rect 34860 44940 34916 44942
rect 34748 44492 34804 44548
rect 34636 44156 34692 44212
rect 34524 42700 34580 42756
rect 34412 42530 34468 42532
rect 34412 42478 34414 42530
rect 34414 42478 34466 42530
rect 34466 42478 34468 42530
rect 34412 42476 34468 42478
rect 34524 42082 34580 42084
rect 34524 42030 34526 42082
rect 34526 42030 34578 42082
rect 34578 42030 34580 42082
rect 34524 42028 34580 42030
rect 33628 41244 33684 41300
rect 29820 40348 29876 40404
rect 30604 40460 30660 40516
rect 32508 39340 32564 39396
rect 30716 39004 30772 39060
rect 29372 38668 29428 38724
rect 33180 40348 33236 40404
rect 34076 41692 34132 41748
rect 33852 41074 33908 41076
rect 33852 41022 33854 41074
rect 33854 41022 33906 41074
rect 33906 41022 33908 41074
rect 33852 41020 33908 41022
rect 33964 40514 34020 40516
rect 33964 40462 33966 40514
rect 33966 40462 34018 40514
rect 34018 40462 34020 40514
rect 33964 40460 34020 40462
rect 34300 41074 34356 41076
rect 34300 41022 34302 41074
rect 34302 41022 34354 41074
rect 34354 41022 34356 41074
rect 34300 41020 34356 41022
rect 34300 40572 34356 40628
rect 33516 39618 33572 39620
rect 33516 39566 33518 39618
rect 33518 39566 33570 39618
rect 33570 39566 33572 39618
rect 33516 39564 33572 39566
rect 34188 39618 34244 39620
rect 34188 39566 34190 39618
rect 34190 39566 34242 39618
rect 34242 39566 34244 39618
rect 34188 39564 34244 39566
rect 33628 39394 33684 39396
rect 33628 39342 33630 39394
rect 33630 39342 33682 39394
rect 33682 39342 33684 39394
rect 33628 39340 33684 39342
rect 29820 38332 29876 38388
rect 29708 38274 29764 38276
rect 29708 38222 29710 38274
rect 29710 38222 29762 38274
rect 29762 38222 29764 38274
rect 29708 38220 29764 38222
rect 29036 37436 29092 37492
rect 29484 38050 29540 38052
rect 29484 37998 29486 38050
rect 29486 37998 29538 38050
rect 29538 37998 29540 38050
rect 29484 37996 29540 37998
rect 30828 37324 30884 37380
rect 30156 36204 30212 36260
rect 29484 35586 29540 35588
rect 29484 35534 29486 35586
rect 29486 35534 29538 35586
rect 29538 35534 29540 35586
rect 29484 35532 29540 35534
rect 29036 34748 29092 34804
rect 29484 34972 29540 35028
rect 27916 32396 27972 32452
rect 27020 31276 27076 31332
rect 28140 31554 28196 31556
rect 28140 31502 28142 31554
rect 28142 31502 28194 31554
rect 28194 31502 28196 31554
rect 28140 31500 28196 31502
rect 27468 31276 27524 31332
rect 26460 30940 26516 30996
rect 25452 30044 25508 30100
rect 26348 29986 26404 29988
rect 26348 29934 26350 29986
rect 26350 29934 26402 29986
rect 26402 29934 26404 29986
rect 26348 29932 26404 29934
rect 27020 29986 27076 29988
rect 27020 29934 27022 29986
rect 27022 29934 27074 29986
rect 27074 29934 27076 29986
rect 27020 29932 27076 29934
rect 25676 28476 25732 28532
rect 26908 29484 26964 29540
rect 25676 27244 25732 27300
rect 26012 28364 26068 28420
rect 27132 28812 27188 28868
rect 26460 28364 26516 28420
rect 26796 28140 26852 28196
rect 25900 26236 25956 26292
rect 25900 25506 25956 25508
rect 25900 25454 25902 25506
rect 25902 25454 25954 25506
rect 25954 25454 25956 25506
rect 25900 25452 25956 25454
rect 26908 27746 26964 27748
rect 26908 27694 26910 27746
rect 26910 27694 26962 27746
rect 26962 27694 26964 27746
rect 26908 27692 26964 27694
rect 27244 27692 27300 27748
rect 27692 30994 27748 30996
rect 27692 30942 27694 30994
rect 27694 30942 27746 30994
rect 27746 30942 27748 30994
rect 27692 30940 27748 30942
rect 28140 30994 28196 30996
rect 28140 30942 28142 30994
rect 28142 30942 28194 30994
rect 28194 30942 28196 30994
rect 28140 30940 28196 30942
rect 27580 30828 27636 30884
rect 28588 32060 28644 32116
rect 27916 29650 27972 29652
rect 27916 29598 27918 29650
rect 27918 29598 27970 29650
rect 27970 29598 27972 29650
rect 27916 29596 27972 29598
rect 27580 28642 27636 28644
rect 27580 28590 27582 28642
rect 27582 28590 27634 28642
rect 27634 28590 27636 28642
rect 27580 28588 27636 28590
rect 27580 27298 27636 27300
rect 27580 27246 27582 27298
rect 27582 27246 27634 27298
rect 27634 27246 27636 27298
rect 27580 27244 27636 27246
rect 27580 26850 27636 26852
rect 27580 26798 27582 26850
rect 27582 26798 27634 26850
rect 27634 26798 27636 26850
rect 27580 26796 27636 26798
rect 27692 26684 27748 26740
rect 27580 26460 27636 26516
rect 28028 29260 28084 29316
rect 28140 28812 28196 28868
rect 28028 28588 28084 28644
rect 27916 28364 27972 28420
rect 27916 28140 27972 28196
rect 28252 28140 28308 28196
rect 28588 31500 28644 31556
rect 29484 31724 29540 31780
rect 29708 34748 29764 34804
rect 29260 31554 29316 31556
rect 29260 31502 29262 31554
rect 29262 31502 29314 31554
rect 29314 31502 29316 31554
rect 29260 31500 29316 31502
rect 29708 31500 29764 31556
rect 29932 34636 29988 34692
rect 29596 31276 29652 31332
rect 28700 30156 28756 30212
rect 29148 30210 29204 30212
rect 29148 30158 29150 30210
rect 29150 30158 29202 30210
rect 29202 30158 29204 30210
rect 29148 30156 29204 30158
rect 29932 31164 29988 31220
rect 29708 30098 29764 30100
rect 29708 30046 29710 30098
rect 29710 30046 29762 30098
rect 29762 30046 29764 30098
rect 29708 30044 29764 30046
rect 29596 29596 29652 29652
rect 28812 29314 28868 29316
rect 28812 29262 28814 29314
rect 28814 29262 28866 29314
rect 28866 29262 28868 29314
rect 28812 29260 28868 29262
rect 28140 26684 28196 26740
rect 28028 26460 28084 26516
rect 25564 25282 25620 25284
rect 25564 25230 25566 25282
rect 25566 25230 25618 25282
rect 25618 25230 25620 25282
rect 25564 25228 25620 25230
rect 25564 24780 25620 24836
rect 27132 25676 27188 25732
rect 26572 25228 26628 25284
rect 26124 24834 26180 24836
rect 26124 24782 26126 24834
rect 26126 24782 26178 24834
rect 26178 24782 26180 24834
rect 26124 24780 26180 24782
rect 26460 25116 26516 25172
rect 26908 25228 26964 25284
rect 27132 25116 27188 25172
rect 26908 24556 26964 24612
rect 26236 23996 26292 24052
rect 26012 22988 26068 23044
rect 26012 22316 26068 22372
rect 25228 20860 25284 20916
rect 27916 25506 27972 25508
rect 27916 25454 27918 25506
rect 27918 25454 27970 25506
rect 27970 25454 27972 25506
rect 27916 25452 27972 25454
rect 27468 24610 27524 24612
rect 27468 24558 27470 24610
rect 27470 24558 27522 24610
rect 27522 24558 27524 24610
rect 27468 24556 27524 24558
rect 27356 23042 27412 23044
rect 27356 22990 27358 23042
rect 27358 22990 27410 23042
rect 27410 22990 27412 23042
rect 27356 22988 27412 22990
rect 28140 25340 28196 25396
rect 28588 28476 28644 28532
rect 28140 24610 28196 24612
rect 28140 24558 28142 24610
rect 28142 24558 28194 24610
rect 28194 24558 28196 24610
rect 28140 24556 28196 24558
rect 27580 22258 27636 22260
rect 27580 22206 27582 22258
rect 27582 22206 27634 22258
rect 27634 22206 27636 22258
rect 27580 22204 27636 22206
rect 26796 20300 26852 20356
rect 26124 20018 26180 20020
rect 26124 19966 26126 20018
rect 26126 19966 26178 20018
rect 26178 19966 26180 20018
rect 26124 19964 26180 19966
rect 26572 20018 26628 20020
rect 26572 19966 26574 20018
rect 26574 19966 26626 20018
rect 26626 19966 26628 20018
rect 26572 19964 26628 19966
rect 26572 19404 26628 19460
rect 25340 19180 25396 19236
rect 25116 18508 25172 18564
rect 24892 18284 24948 18340
rect 26236 18396 26292 18452
rect 26572 18508 26628 18564
rect 24444 15932 24500 15988
rect 24668 17500 24724 17556
rect 24892 16716 24948 16772
rect 25788 17554 25844 17556
rect 25788 17502 25790 17554
rect 25790 17502 25842 17554
rect 25842 17502 25844 17554
rect 25788 17500 25844 17502
rect 25228 16716 25284 16772
rect 25116 16098 25172 16100
rect 25116 16046 25118 16098
rect 25118 16046 25170 16098
rect 25170 16046 25172 16098
rect 25116 16044 25172 16046
rect 25676 17442 25732 17444
rect 25676 17390 25678 17442
rect 25678 17390 25730 17442
rect 25730 17390 25732 17442
rect 25676 17388 25732 17390
rect 24108 15260 24164 15316
rect 23436 13356 23492 13412
rect 23548 12290 23604 12292
rect 23548 12238 23550 12290
rect 23550 12238 23602 12290
rect 23602 12238 23604 12290
rect 23548 12236 23604 12238
rect 20860 8540 20916 8596
rect 21756 9212 21812 9268
rect 21756 8316 21812 8372
rect 16268 7308 16324 7364
rect 14812 6748 14868 6804
rect 16380 6802 16436 6804
rect 16380 6750 16382 6802
rect 16382 6750 16434 6802
rect 16434 6750 16436 6802
rect 16380 6748 16436 6750
rect 17052 7308 17108 7364
rect 19516 8034 19572 8036
rect 19516 7982 19518 8034
rect 19518 7982 19570 8034
rect 19570 7982 19572 8034
rect 19516 7980 19572 7982
rect 18508 7586 18564 7588
rect 18508 7534 18510 7586
rect 18510 7534 18562 7586
rect 18562 7534 18564 7586
rect 18508 7532 18564 7534
rect 20636 8258 20692 8260
rect 20636 8206 20638 8258
rect 20638 8206 20690 8258
rect 20690 8206 20692 8258
rect 20636 8204 20692 8206
rect 20300 7980 20356 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19180 7532 19236 7588
rect 23436 10722 23492 10724
rect 23436 10670 23438 10722
rect 23438 10670 23490 10722
rect 23490 10670 23492 10722
rect 23436 10668 23492 10670
rect 24332 14530 24388 14532
rect 24332 14478 24334 14530
rect 24334 14478 24386 14530
rect 24386 14478 24388 14530
rect 24332 14476 24388 14478
rect 24668 14476 24724 14532
rect 24220 14306 24276 14308
rect 24220 14254 24222 14306
rect 24222 14254 24274 14306
rect 24274 14254 24276 14306
rect 24220 14252 24276 14254
rect 24668 13746 24724 13748
rect 24668 13694 24670 13746
rect 24670 13694 24722 13746
rect 24722 13694 24724 13746
rect 24668 13692 24724 13694
rect 24220 13580 24276 13636
rect 24444 13580 24500 13636
rect 24444 12236 24500 12292
rect 23772 12178 23828 12180
rect 23772 12126 23774 12178
rect 23774 12126 23826 12178
rect 23826 12126 23828 12178
rect 23772 12124 23828 12126
rect 24332 12178 24388 12180
rect 24332 12126 24334 12178
rect 24334 12126 24386 12178
rect 24386 12126 24388 12178
rect 24332 12124 24388 12126
rect 23996 12012 24052 12068
rect 23772 11900 23828 11956
rect 23772 10556 23828 10612
rect 23436 9154 23492 9156
rect 23436 9102 23438 9154
rect 23438 9102 23490 9154
rect 23490 9102 23492 9154
rect 23436 9100 23492 9102
rect 22652 7980 22708 8036
rect 22540 7644 22596 7700
rect 22316 7532 22372 7588
rect 18732 7474 18788 7476
rect 18732 7422 18734 7474
rect 18734 7422 18786 7474
rect 18786 7422 18788 7474
rect 18732 7420 18788 7422
rect 17948 7308 18004 7364
rect 17724 7196 17780 7252
rect 18396 7250 18452 7252
rect 18396 7198 18398 7250
rect 18398 7198 18450 7250
rect 18450 7198 18452 7250
rect 18396 7196 18452 7198
rect 19292 7362 19348 7364
rect 19292 7310 19294 7362
rect 19294 7310 19346 7362
rect 19346 7310 19348 7362
rect 19292 7308 19348 7310
rect 18396 5180 18452 5236
rect 16716 5122 16772 5124
rect 16716 5070 16718 5122
rect 16718 5070 16770 5122
rect 16770 5070 16772 5122
rect 16716 5068 16772 5070
rect 14364 4508 14420 4564
rect 14924 4562 14980 4564
rect 14924 4510 14926 4562
rect 14926 4510 14978 4562
rect 14978 4510 14980 4562
rect 14924 4508 14980 4510
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 7196 3388 7252 3444
rect 10108 3442 10164 3444
rect 10108 3390 10110 3442
rect 10110 3390 10162 3442
rect 10162 3390 10164 3442
rect 10108 3388 10164 3390
rect 18844 5234 18900 5236
rect 18844 5182 18846 5234
rect 18846 5182 18898 5234
rect 18898 5182 18900 5234
rect 18844 5180 18900 5182
rect 19180 5068 19236 5124
rect 19516 5740 19572 5796
rect 19292 4898 19348 4900
rect 19292 4846 19294 4898
rect 19294 4846 19346 4898
rect 19346 4846 19348 4898
rect 19292 4844 19348 4846
rect 19852 6860 19908 6916
rect 22316 6860 22372 6916
rect 22204 6748 22260 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 22988 8204 23044 8260
rect 23212 8092 23268 8148
rect 23100 8034 23156 8036
rect 23100 7982 23102 8034
rect 23102 7982 23154 8034
rect 23154 7982 23156 8034
rect 23100 7980 23156 7982
rect 23100 7698 23156 7700
rect 23100 7646 23102 7698
rect 23102 7646 23154 7698
rect 23154 7646 23156 7698
rect 23100 7644 23156 7646
rect 23324 7756 23380 7812
rect 23548 8146 23604 8148
rect 23548 8094 23550 8146
rect 23550 8094 23602 8146
rect 23602 8094 23604 8146
rect 23548 8092 23604 8094
rect 23436 7532 23492 7588
rect 23212 7474 23268 7476
rect 23212 7422 23214 7474
rect 23214 7422 23266 7474
rect 23266 7422 23268 7474
rect 23212 7420 23268 7422
rect 22988 6748 23044 6804
rect 22988 6076 23044 6132
rect 22540 6018 22596 6020
rect 22540 5966 22542 6018
rect 22542 5966 22594 6018
rect 22594 5966 22596 6018
rect 22540 5964 22596 5966
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21644 5122 21700 5124
rect 21644 5070 21646 5122
rect 21646 5070 21698 5122
rect 21698 5070 21700 5122
rect 21644 5068 21700 5070
rect 22428 5794 22484 5796
rect 22428 5742 22430 5794
rect 22430 5742 22482 5794
rect 22482 5742 22484 5794
rect 22428 5740 22484 5742
rect 22876 5964 22932 6020
rect 22652 5180 22708 5236
rect 22428 5068 22484 5124
rect 23772 7532 23828 7588
rect 24220 10722 24276 10724
rect 24220 10670 24222 10722
rect 24222 10670 24274 10722
rect 24274 10670 24276 10722
rect 24220 10668 24276 10670
rect 24668 12178 24724 12180
rect 24668 12126 24670 12178
rect 24670 12126 24722 12178
rect 24722 12126 24724 12178
rect 24668 12124 24724 12126
rect 25340 15708 25396 15764
rect 26012 14530 26068 14532
rect 26012 14478 26014 14530
rect 26014 14478 26066 14530
rect 26066 14478 26068 14530
rect 26012 14476 26068 14478
rect 25340 14252 25396 14308
rect 26124 14306 26180 14308
rect 26124 14254 26126 14306
rect 26126 14254 26178 14306
rect 26178 14254 26180 14306
rect 26124 14252 26180 14254
rect 25340 13634 25396 13636
rect 25340 13582 25342 13634
rect 25342 13582 25394 13634
rect 25394 13582 25396 13634
rect 25340 13580 25396 13582
rect 25788 13580 25844 13636
rect 26124 13634 26180 13636
rect 26124 13582 26126 13634
rect 26126 13582 26178 13634
rect 26178 13582 26180 13634
rect 26124 13580 26180 13582
rect 25228 11900 25284 11956
rect 26124 12796 26180 12852
rect 25788 11788 25844 11844
rect 25900 12124 25956 12180
rect 26124 11788 26180 11844
rect 26348 11228 26404 11284
rect 25228 10722 25284 10724
rect 25228 10670 25230 10722
rect 25230 10670 25282 10722
rect 25282 10670 25284 10722
rect 25228 10668 25284 10670
rect 26236 10220 26292 10276
rect 26012 10108 26068 10164
rect 27132 18562 27188 18564
rect 27132 18510 27134 18562
rect 27134 18510 27186 18562
rect 27186 18510 27188 18562
rect 27132 18508 27188 18510
rect 27020 18450 27076 18452
rect 27020 18398 27022 18450
rect 27022 18398 27074 18450
rect 27074 18398 27076 18450
rect 27020 18396 27076 18398
rect 27580 18956 27636 19012
rect 30156 35532 30212 35588
rect 30156 35026 30212 35028
rect 30156 34974 30158 35026
rect 30158 34974 30210 35026
rect 30210 34974 30212 35026
rect 30156 34972 30212 34974
rect 30044 28476 30100 28532
rect 30268 30044 30324 30100
rect 29708 28140 29764 28196
rect 29036 26908 29092 26964
rect 28588 26124 28644 26180
rect 28924 26572 28980 26628
rect 28476 25282 28532 25284
rect 28476 25230 28478 25282
rect 28478 25230 28530 25282
rect 28530 25230 28532 25282
rect 28476 25228 28532 25230
rect 28588 24892 28644 24948
rect 28364 24834 28420 24836
rect 28364 24782 28366 24834
rect 28366 24782 28418 24834
rect 28418 24782 28420 24834
rect 28364 24780 28420 24782
rect 29148 26796 29204 26852
rect 30604 34860 30660 34916
rect 30604 34690 30660 34692
rect 30604 34638 30606 34690
rect 30606 34638 30658 34690
rect 30658 34638 30660 34690
rect 30604 34636 30660 34638
rect 30604 34018 30660 34020
rect 30604 33966 30606 34018
rect 30606 33966 30658 34018
rect 30658 33966 30660 34018
rect 30604 33964 30660 33966
rect 31836 36316 31892 36372
rect 31612 35698 31668 35700
rect 31612 35646 31614 35698
rect 31614 35646 31666 35698
rect 31666 35646 31668 35698
rect 31612 35644 31668 35646
rect 31052 34972 31108 35028
rect 32620 35922 32676 35924
rect 32620 35870 32622 35922
rect 32622 35870 32674 35922
rect 32674 35870 32676 35922
rect 32620 35868 32676 35870
rect 32284 35644 32340 35700
rect 31276 34860 31332 34916
rect 30940 34748 30996 34804
rect 31948 34748 32004 34804
rect 30828 32284 30884 32340
rect 31164 33068 31220 33124
rect 32396 34860 32452 34916
rect 33516 38108 33572 38164
rect 33180 35698 33236 35700
rect 33180 35646 33182 35698
rect 33182 35646 33234 35698
rect 33234 35646 33236 35698
rect 33180 35644 33236 35646
rect 33516 35084 33572 35140
rect 33404 34860 33460 34916
rect 32620 34636 32676 34692
rect 33292 34242 33348 34244
rect 33292 34190 33294 34242
rect 33294 34190 33346 34242
rect 33346 34190 33348 34242
rect 33292 34188 33348 34190
rect 32396 33964 32452 34020
rect 32396 33404 32452 33460
rect 32844 33458 32900 33460
rect 32844 33406 32846 33458
rect 32846 33406 32898 33458
rect 32898 33406 32900 33458
rect 32844 33404 32900 33406
rect 31164 31948 31220 32004
rect 30492 31388 30548 31444
rect 30604 29708 30660 29764
rect 30828 30828 30884 30884
rect 31724 31724 31780 31780
rect 32284 31778 32340 31780
rect 32284 31726 32286 31778
rect 32286 31726 32338 31778
rect 32338 31726 32340 31778
rect 32284 31724 32340 31726
rect 31612 31388 31668 31444
rect 31276 30940 31332 30996
rect 31388 30210 31444 30212
rect 31388 30158 31390 30210
rect 31390 30158 31442 30210
rect 31442 30158 31444 30210
rect 31388 30156 31444 30158
rect 31276 29986 31332 29988
rect 31276 29934 31278 29986
rect 31278 29934 31330 29986
rect 31330 29934 31332 29986
rect 31276 29932 31332 29934
rect 30492 28418 30548 28420
rect 30492 28366 30494 28418
rect 30494 28366 30546 28418
rect 30546 28366 30548 28418
rect 30492 28364 30548 28366
rect 30828 29372 30884 29428
rect 31612 30156 31668 30212
rect 31948 29986 32004 29988
rect 31948 29934 31950 29986
rect 31950 29934 32002 29986
rect 32002 29934 32004 29986
rect 31948 29932 32004 29934
rect 30268 26348 30324 26404
rect 30380 27916 30436 27972
rect 29820 26124 29876 26180
rect 30268 26178 30324 26180
rect 30268 26126 30270 26178
rect 30270 26126 30322 26178
rect 30322 26126 30324 26178
rect 30268 26124 30324 26126
rect 29372 25506 29428 25508
rect 29372 25454 29374 25506
rect 29374 25454 29426 25506
rect 29426 25454 29428 25506
rect 29372 25452 29428 25454
rect 29932 25394 29988 25396
rect 29932 25342 29934 25394
rect 29934 25342 29986 25394
rect 29986 25342 29988 25394
rect 29932 25340 29988 25342
rect 28924 24780 28980 24836
rect 29708 24834 29764 24836
rect 29708 24782 29710 24834
rect 29710 24782 29762 24834
rect 29762 24782 29764 24834
rect 29708 24780 29764 24782
rect 29036 24722 29092 24724
rect 29036 24670 29038 24722
rect 29038 24670 29090 24722
rect 29090 24670 29092 24722
rect 29036 24668 29092 24670
rect 28588 22988 28644 23044
rect 29260 22652 29316 22708
rect 29148 22428 29204 22484
rect 30828 28364 30884 28420
rect 30716 27132 30772 27188
rect 30604 26962 30660 26964
rect 30604 26910 30606 26962
rect 30606 26910 30658 26962
rect 30658 26910 30660 26962
rect 30604 26908 30660 26910
rect 31388 28700 31444 28756
rect 31276 27970 31332 27972
rect 31276 27918 31278 27970
rect 31278 27918 31330 27970
rect 31330 27918 31332 27970
rect 31276 27916 31332 27918
rect 31724 29708 31780 29764
rect 32172 29426 32228 29428
rect 32172 29374 32174 29426
rect 32174 29374 32226 29426
rect 32226 29374 32228 29426
rect 32172 29372 32228 29374
rect 31052 27244 31108 27300
rect 31724 28476 31780 28532
rect 31612 26908 31668 26964
rect 30828 26236 30884 26292
rect 30492 25452 30548 25508
rect 30268 24946 30324 24948
rect 30268 24894 30270 24946
rect 30270 24894 30322 24946
rect 30322 24894 30324 24946
rect 30268 24892 30324 24894
rect 30604 24780 30660 24836
rect 29484 22092 29540 22148
rect 30044 21644 30100 21700
rect 29148 20690 29204 20692
rect 29148 20638 29150 20690
rect 29150 20638 29202 20690
rect 29202 20638 29204 20690
rect 29148 20636 29204 20638
rect 29932 20914 29988 20916
rect 29932 20862 29934 20914
rect 29934 20862 29986 20914
rect 29986 20862 29988 20914
rect 29932 20860 29988 20862
rect 30380 22146 30436 22148
rect 30380 22094 30382 22146
rect 30382 22094 30434 22146
rect 30434 22094 30436 22146
rect 30380 22092 30436 22094
rect 31836 27244 31892 27300
rect 32284 27186 32340 27188
rect 32284 27134 32286 27186
rect 32286 27134 32338 27186
rect 32338 27134 32340 27186
rect 32284 27132 32340 27134
rect 31948 27020 32004 27076
rect 31164 25676 31220 25732
rect 31276 26124 31332 26180
rect 31724 25564 31780 25620
rect 31276 25228 31332 25284
rect 30828 22092 30884 22148
rect 31052 24892 31108 24948
rect 30380 21420 30436 21476
rect 31164 22428 31220 22484
rect 30044 20636 30100 20692
rect 29484 19852 29540 19908
rect 30828 20690 30884 20692
rect 30828 20638 30830 20690
rect 30830 20638 30882 20690
rect 30882 20638 30884 20690
rect 30828 20636 30884 20638
rect 30268 20018 30324 20020
rect 30268 19966 30270 20018
rect 30270 19966 30322 20018
rect 30322 19966 30324 20018
rect 30268 19964 30324 19966
rect 29372 19234 29428 19236
rect 29372 19182 29374 19234
rect 29374 19182 29426 19234
rect 29426 19182 29428 19234
rect 29372 19180 29428 19182
rect 28476 19068 28532 19124
rect 29036 19010 29092 19012
rect 29036 18958 29038 19010
rect 29038 18958 29090 19010
rect 29090 18958 29092 19010
rect 29036 18956 29092 18958
rect 29260 19010 29316 19012
rect 29260 18958 29262 19010
rect 29262 18958 29314 19010
rect 29314 18958 29316 19010
rect 29260 18956 29316 18958
rect 28252 17388 28308 17444
rect 28812 15932 28868 15988
rect 29260 15708 29316 15764
rect 30268 19234 30324 19236
rect 30268 19182 30270 19234
rect 30270 19182 30322 19234
rect 30322 19182 30324 19234
rect 30268 19180 30324 19182
rect 29820 19010 29876 19012
rect 29820 18958 29822 19010
rect 29822 18958 29874 19010
rect 29874 18958 29876 19010
rect 29820 18956 29876 18958
rect 30492 19740 30548 19796
rect 30828 19964 30884 20020
rect 29932 18284 29988 18340
rect 30268 17052 30324 17108
rect 28476 15314 28532 15316
rect 28476 15262 28478 15314
rect 28478 15262 28530 15314
rect 28530 15262 28532 15314
rect 28476 15260 28532 15262
rect 26796 14924 26852 14980
rect 26572 13746 26628 13748
rect 26572 13694 26574 13746
rect 26574 13694 26626 13746
rect 26626 13694 26628 13746
rect 26572 13692 26628 13694
rect 26684 13244 26740 13300
rect 26572 12738 26628 12740
rect 26572 12686 26574 12738
rect 26574 12686 26626 12738
rect 26626 12686 26628 12738
rect 26572 12684 26628 12686
rect 26684 11788 26740 11844
rect 27020 13244 27076 13300
rect 27132 12796 27188 12852
rect 27132 12348 27188 12404
rect 26908 12066 26964 12068
rect 26908 12014 26910 12066
rect 26910 12014 26962 12066
rect 26962 12014 26964 12066
rect 26908 12012 26964 12014
rect 26796 11282 26852 11284
rect 26796 11230 26798 11282
rect 26798 11230 26850 11282
rect 26850 11230 26852 11282
rect 26796 11228 26852 11230
rect 25340 8540 25396 8596
rect 26236 8370 26292 8372
rect 26236 8318 26238 8370
rect 26238 8318 26290 8370
rect 26290 8318 26292 8370
rect 26236 8316 26292 8318
rect 24556 8092 24612 8148
rect 25452 8092 25508 8148
rect 24780 7980 24836 8036
rect 25004 7756 25060 7812
rect 23884 6748 23940 6804
rect 23660 6076 23716 6132
rect 24220 6466 24276 6468
rect 24220 6414 24222 6466
rect 24222 6414 24274 6466
rect 24274 6414 24276 6466
rect 24220 6412 24276 6414
rect 24220 6130 24276 6132
rect 24220 6078 24222 6130
rect 24222 6078 24274 6130
rect 24274 6078 24276 6130
rect 24220 6076 24276 6078
rect 24444 6130 24500 6132
rect 24444 6078 24446 6130
rect 24446 6078 24498 6130
rect 24498 6078 24500 6130
rect 24444 6076 24500 6078
rect 26012 8092 26068 8148
rect 26348 8034 26404 8036
rect 26348 7982 26350 8034
rect 26350 7982 26402 8034
rect 26402 7982 26404 8034
rect 26348 7980 26404 7982
rect 25900 7756 25956 7812
rect 26236 7474 26292 7476
rect 26236 7422 26238 7474
rect 26238 7422 26290 7474
rect 26290 7422 26292 7474
rect 26236 7420 26292 7422
rect 25452 6972 25508 7028
rect 27580 14924 27636 14980
rect 27356 13634 27412 13636
rect 27356 13582 27358 13634
rect 27358 13582 27410 13634
rect 27410 13582 27412 13634
rect 27356 13580 27412 13582
rect 28252 12402 28308 12404
rect 28252 12350 28254 12402
rect 28254 12350 28306 12402
rect 28306 12350 28308 12402
rect 28252 12348 28308 12350
rect 27020 11394 27076 11396
rect 27020 11342 27022 11394
rect 27022 11342 27074 11394
rect 27074 11342 27076 11394
rect 27020 11340 27076 11342
rect 27132 10220 27188 10276
rect 27132 9826 27188 9828
rect 27132 9774 27134 9826
rect 27134 9774 27186 9826
rect 27186 9774 27188 9826
rect 27132 9772 27188 9774
rect 27244 8370 27300 8372
rect 27244 8318 27246 8370
rect 27246 8318 27298 8370
rect 27298 8318 27300 8370
rect 27244 8316 27300 8318
rect 27020 7308 27076 7364
rect 27020 6972 27076 7028
rect 26684 6076 26740 6132
rect 24556 5906 24612 5908
rect 24556 5854 24558 5906
rect 24558 5854 24610 5906
rect 24610 5854 24612 5906
rect 24556 5852 24612 5854
rect 21420 4898 21476 4900
rect 21420 4846 21422 4898
rect 21422 4846 21474 4898
rect 21474 4846 21476 4898
rect 21420 4844 21476 4846
rect 23548 5180 23604 5236
rect 18396 3612 18452 3668
rect 11900 3388 11956 3444
rect 12460 3442 12516 3444
rect 12460 3390 12462 3442
rect 12462 3390 12514 3442
rect 12514 3390 12516 3442
rect 12460 3388 12516 3390
rect 25340 5122 25396 5124
rect 25340 5070 25342 5122
rect 25342 5070 25394 5122
rect 25394 5070 25396 5122
rect 25340 5068 25396 5070
rect 24668 3554 24724 3556
rect 24668 3502 24670 3554
rect 24670 3502 24722 3554
rect 24722 3502 24724 3554
rect 24668 3500 24724 3502
rect 23548 3388 23604 3444
rect 16156 3276 16212 3332
rect 16940 3330 16996 3332
rect 16940 3278 16942 3330
rect 16942 3278 16994 3330
rect 16994 3278 16996 3330
rect 16940 3276 16996 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25788 5122 25844 5124
rect 25788 5070 25790 5122
rect 25790 5070 25842 5122
rect 25842 5070 25844 5122
rect 25788 5068 25844 5070
rect 26908 5068 26964 5124
rect 27244 5852 27300 5908
rect 29596 15314 29652 15316
rect 29596 15262 29598 15314
rect 29598 15262 29650 15314
rect 29650 15262 29652 15314
rect 29596 15260 29652 15262
rect 29484 14812 29540 14868
rect 29484 14252 29540 14308
rect 30156 14588 30212 14644
rect 29372 13244 29428 13300
rect 30156 13132 30212 13188
rect 30716 14252 30772 14308
rect 30268 12348 30324 12404
rect 30716 12012 30772 12068
rect 29484 11564 29540 11620
rect 29260 11394 29316 11396
rect 29260 11342 29262 11394
rect 29262 11342 29314 11394
rect 29314 11342 29316 11394
rect 29260 11340 29316 11342
rect 30380 10892 30436 10948
rect 30156 10780 30212 10836
rect 29932 10556 29988 10612
rect 29148 9772 29204 9828
rect 29484 10108 29540 10164
rect 32172 25676 32228 25732
rect 31948 25618 32004 25620
rect 31948 25566 31950 25618
rect 31950 25566 32002 25618
rect 32002 25566 32004 25618
rect 31948 25564 32004 25566
rect 32060 24780 32116 24836
rect 34636 35586 34692 35588
rect 34636 35534 34638 35586
rect 34638 35534 34690 35586
rect 34690 35534 34692 35586
rect 34636 35532 34692 35534
rect 34076 35308 34132 35364
rect 34636 35308 34692 35364
rect 37324 47234 37380 47236
rect 37324 47182 37326 47234
rect 37326 47182 37378 47234
rect 37378 47182 37380 47234
rect 37324 47180 37380 47182
rect 36876 46674 36932 46676
rect 36876 46622 36878 46674
rect 36878 46622 36930 46674
rect 36930 46622 36932 46674
rect 36876 46620 36932 46622
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35980 45724 36036 45780
rect 35308 45052 35364 45108
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35532 44546 35588 44548
rect 35532 44494 35534 44546
rect 35534 44494 35586 44546
rect 35586 44494 35588 44546
rect 35532 44492 35588 44494
rect 35084 44434 35140 44436
rect 35084 44382 35086 44434
rect 35086 44382 35138 44434
rect 35138 44382 35140 44434
rect 35084 44380 35140 44382
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35084 42588 35140 42644
rect 35084 42082 35140 42084
rect 35084 42030 35086 42082
rect 35086 42030 35138 42082
rect 35138 42030 35140 42082
rect 35084 42028 35140 42030
rect 34972 41746 35028 41748
rect 34972 41694 34974 41746
rect 34974 41694 35026 41746
rect 35026 41694 35028 41746
rect 34972 41692 35028 41694
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35756 44210 35812 44212
rect 35756 44158 35758 44210
rect 35758 44158 35810 44210
rect 35810 44158 35812 44210
rect 35756 44156 35812 44158
rect 36092 45052 36148 45108
rect 36092 43932 36148 43988
rect 35980 43426 36036 43428
rect 35980 43374 35982 43426
rect 35982 43374 36034 43426
rect 36034 43374 36036 43426
rect 35980 43372 36036 43374
rect 36428 46172 36484 46228
rect 41132 49922 41188 49924
rect 41132 49870 41134 49922
rect 41134 49870 41186 49922
rect 41186 49870 41188 49922
rect 41132 49868 41188 49870
rect 39900 49698 39956 49700
rect 39900 49646 39902 49698
rect 39902 49646 39954 49698
rect 39954 49646 39956 49698
rect 39900 49644 39956 49646
rect 39788 48860 39844 48916
rect 39228 47628 39284 47684
rect 37660 46172 37716 46228
rect 37324 45724 37380 45780
rect 37884 45724 37940 45780
rect 37100 45052 37156 45108
rect 38220 45106 38276 45108
rect 38220 45054 38222 45106
rect 38222 45054 38274 45106
rect 38274 45054 38276 45106
rect 38220 45052 38276 45054
rect 37212 44940 37268 44996
rect 37100 44380 37156 44436
rect 37772 44156 37828 44212
rect 36316 43708 36372 43764
rect 39228 47180 39284 47236
rect 38892 46284 38948 46340
rect 38780 45052 38836 45108
rect 38556 44322 38612 44324
rect 38556 44270 38558 44322
rect 38558 44270 38610 44322
rect 38610 44270 38612 44322
rect 38556 44268 38612 44270
rect 39004 44322 39060 44324
rect 39004 44270 39006 44322
rect 39006 44270 39058 44322
rect 39058 44270 39060 44322
rect 39004 44268 39060 44270
rect 37884 43820 37940 43876
rect 38780 43932 38836 43988
rect 40908 49698 40964 49700
rect 40908 49646 40910 49698
rect 40910 49646 40962 49698
rect 40962 49646 40964 49698
rect 40908 49644 40964 49646
rect 40236 47404 40292 47460
rect 41132 48860 41188 48916
rect 40012 46956 40068 47012
rect 39900 46620 39956 46676
rect 39452 44268 39508 44324
rect 39452 43708 39508 43764
rect 35980 42642 36036 42644
rect 35980 42590 35982 42642
rect 35982 42590 36034 42642
rect 36034 42590 36036 42642
rect 35980 42588 36036 42590
rect 35868 42476 35924 42532
rect 38556 42754 38612 42756
rect 38556 42702 38558 42754
rect 38558 42702 38610 42754
rect 38610 42702 38612 42754
rect 38556 42700 38612 42702
rect 35868 42028 35924 42084
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 38220 42530 38276 42532
rect 38220 42478 38222 42530
rect 38222 42478 38274 42530
rect 38274 42478 38276 42530
rect 38220 42476 38276 42478
rect 36204 41132 36260 41188
rect 36988 42252 37044 42308
rect 36652 40908 36708 40964
rect 37100 41916 37156 41972
rect 38108 41244 38164 41300
rect 37212 41186 37268 41188
rect 37212 41134 37214 41186
rect 37214 41134 37266 41186
rect 37266 41134 37268 41186
rect 37212 41132 37268 41134
rect 38556 41298 38612 41300
rect 38556 41246 38558 41298
rect 38558 41246 38610 41298
rect 38610 41246 38612 41298
rect 38556 41244 38612 41246
rect 37100 41020 37156 41076
rect 37324 40962 37380 40964
rect 37324 40910 37326 40962
rect 37326 40910 37378 40962
rect 37378 40910 37380 40962
rect 37324 40908 37380 40910
rect 38556 40684 38612 40740
rect 39452 40684 39508 40740
rect 37996 40236 38052 40292
rect 38780 40290 38836 40292
rect 38780 40238 38782 40290
rect 38782 40238 38834 40290
rect 38834 40238 38836 40290
rect 38780 40236 38836 40238
rect 36988 39788 37044 39844
rect 38780 39116 38836 39172
rect 38108 38780 38164 38836
rect 35532 38108 35588 38164
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 37212 38668 37268 38724
rect 35532 35644 35588 35700
rect 33516 33852 33572 33908
rect 34300 34748 34356 34804
rect 34188 34300 34244 34356
rect 34524 34412 34580 34468
rect 33964 34242 34020 34244
rect 33964 34190 33966 34242
rect 33966 34190 34018 34242
rect 34018 34190 34020 34242
rect 33964 34188 34020 34190
rect 34524 34130 34580 34132
rect 34524 34078 34526 34130
rect 34526 34078 34578 34130
rect 34578 34078 34580 34130
rect 34524 34076 34580 34078
rect 34412 33852 34468 33908
rect 33740 33516 33796 33572
rect 33964 33404 34020 33460
rect 33516 32786 33572 32788
rect 33516 32734 33518 32786
rect 33518 32734 33570 32786
rect 33570 32734 33572 32786
rect 33516 32732 33572 32734
rect 33068 30828 33124 30884
rect 32396 24780 32452 24836
rect 32508 29932 32564 29988
rect 31500 22652 31556 22708
rect 32396 20860 32452 20916
rect 31500 20578 31556 20580
rect 31500 20526 31502 20578
rect 31502 20526 31554 20578
rect 31554 20526 31556 20578
rect 31500 20524 31556 20526
rect 32060 20524 32116 20580
rect 31836 20130 31892 20132
rect 31836 20078 31838 20130
rect 31838 20078 31890 20130
rect 31890 20078 31892 20130
rect 31836 20076 31892 20078
rect 32172 20018 32228 20020
rect 32172 19966 32174 20018
rect 32174 19966 32226 20018
rect 32226 19966 32228 20018
rect 32172 19964 32228 19966
rect 31388 19740 31444 19796
rect 35196 35420 35252 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35532 34802 35588 34804
rect 35532 34750 35534 34802
rect 35534 34750 35586 34802
rect 35586 34750 35588 34802
rect 35532 34748 35588 34750
rect 34860 34300 34916 34356
rect 34636 31948 34692 32004
rect 34972 34188 35028 34244
rect 34300 31106 34356 31108
rect 34300 31054 34302 31106
rect 34302 31054 34354 31106
rect 34354 31054 34356 31106
rect 34300 31052 34356 31054
rect 33740 29820 33796 29876
rect 34188 30156 34244 30212
rect 34076 29708 34132 29764
rect 33516 29484 33572 29540
rect 32732 28476 32788 28532
rect 33516 28252 33572 28308
rect 33628 28700 33684 28756
rect 32732 27356 32788 27412
rect 35196 34300 35252 34356
rect 35420 34412 35476 34468
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35756 34188 35812 34244
rect 35980 38444 36036 38500
rect 36092 35420 36148 35476
rect 35980 35084 36036 35140
rect 37100 38162 37156 38164
rect 37100 38110 37102 38162
rect 37102 38110 37154 38162
rect 37154 38110 37156 38162
rect 37100 38108 37156 38110
rect 38220 38722 38276 38724
rect 38220 38670 38222 38722
rect 38222 38670 38274 38722
rect 38274 38670 38276 38722
rect 38220 38668 38276 38670
rect 39340 39116 39396 39172
rect 38556 38108 38612 38164
rect 37212 34412 37268 34468
rect 35980 34300 36036 34356
rect 35868 34076 35924 34132
rect 35644 33404 35700 33460
rect 35644 32284 35700 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31500 35588 31556
rect 35308 31106 35364 31108
rect 35308 31054 35310 31106
rect 35310 31054 35362 31106
rect 35362 31054 35364 31106
rect 35308 31052 35364 31054
rect 35532 31052 35588 31108
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34860 29932 34916 29988
rect 34300 29372 34356 29428
rect 33628 25228 33684 25284
rect 33964 27804 34020 27860
rect 32620 24556 32676 24612
rect 32732 21308 32788 21364
rect 31276 18844 31332 18900
rect 31836 18844 31892 18900
rect 31500 18620 31556 18676
rect 31500 18450 31556 18452
rect 31500 18398 31502 18450
rect 31502 18398 31554 18450
rect 31554 18398 31556 18450
rect 31500 18396 31556 18398
rect 31612 18338 31668 18340
rect 31612 18286 31614 18338
rect 31614 18286 31666 18338
rect 31666 18286 31668 18338
rect 31612 18284 31668 18286
rect 33964 20972 34020 21028
rect 32956 20914 33012 20916
rect 32956 20862 32958 20914
rect 32958 20862 33010 20914
rect 33010 20862 33012 20914
rect 32956 20860 33012 20862
rect 33516 20524 33572 20580
rect 33180 20130 33236 20132
rect 33180 20078 33182 20130
rect 33182 20078 33234 20130
rect 33234 20078 33236 20130
rect 33180 20076 33236 20078
rect 33068 19964 33124 20020
rect 32732 19292 32788 19348
rect 32844 19628 32900 19684
rect 31948 18562 32004 18564
rect 31948 18510 31950 18562
rect 31950 18510 32002 18562
rect 32002 18510 32004 18562
rect 31948 18508 32004 18510
rect 32172 18450 32228 18452
rect 32172 18398 32174 18450
rect 32174 18398 32226 18450
rect 32226 18398 32228 18450
rect 32172 18396 32228 18398
rect 31836 17948 31892 18004
rect 31724 17836 31780 17892
rect 32508 19180 32564 19236
rect 33628 19234 33684 19236
rect 33628 19182 33630 19234
rect 33630 19182 33682 19234
rect 33682 19182 33684 19234
rect 33628 19180 33684 19182
rect 33404 19068 33460 19124
rect 33740 18844 33796 18900
rect 32508 18562 32564 18564
rect 32508 18510 32510 18562
rect 32510 18510 32562 18562
rect 32562 18510 32564 18562
rect 32508 18508 32564 18510
rect 32620 17890 32676 17892
rect 32620 17838 32622 17890
rect 32622 17838 32674 17890
rect 32674 17838 32676 17890
rect 32620 17836 32676 17838
rect 33180 17724 33236 17780
rect 32396 17612 32452 17668
rect 33068 17612 33124 17668
rect 35084 29596 35140 29652
rect 34972 29538 35028 29540
rect 34972 29486 34974 29538
rect 34974 29486 35026 29538
rect 35026 29486 35028 29538
rect 34972 29484 35028 29486
rect 34524 28140 34580 28196
rect 35644 29932 35700 29988
rect 35532 29538 35588 29540
rect 35532 29486 35534 29538
rect 35534 29486 35586 29538
rect 35586 29486 35588 29538
rect 35532 29484 35588 29486
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34972 28754 35028 28756
rect 34972 28702 34974 28754
rect 34974 28702 35026 28754
rect 35026 28702 35028 28754
rect 34972 28700 35028 28702
rect 35196 28140 35252 28196
rect 34972 28082 35028 28084
rect 34972 28030 34974 28082
rect 34974 28030 35026 28082
rect 35026 28030 35028 28082
rect 34972 28028 35028 28030
rect 34748 27804 34804 27860
rect 34188 27356 34244 27412
rect 34524 27074 34580 27076
rect 34524 27022 34526 27074
rect 34526 27022 34578 27074
rect 34578 27022 34580 27074
rect 34524 27020 34580 27022
rect 37100 33180 37156 33236
rect 36988 32786 37044 32788
rect 36988 32734 36990 32786
rect 36990 32734 37042 32786
rect 37042 32734 37044 32786
rect 36988 32732 37044 32734
rect 37212 33122 37268 33124
rect 37212 33070 37214 33122
rect 37214 33070 37266 33122
rect 37266 33070 37268 33122
rect 37212 33068 37268 33070
rect 36876 29932 36932 29988
rect 35868 29820 35924 29876
rect 35980 29596 36036 29652
rect 35532 28140 35588 28196
rect 35644 27804 35700 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35644 27074 35700 27076
rect 35644 27022 35646 27074
rect 35646 27022 35698 27074
rect 35698 27022 35700 27074
rect 35644 27020 35700 27022
rect 34412 26908 34468 26964
rect 35980 28082 36036 28084
rect 35980 28030 35982 28082
rect 35982 28030 36034 28082
rect 36034 28030 36036 28082
rect 35980 28028 36036 28030
rect 36652 28700 36708 28756
rect 39228 36876 39284 36932
rect 39116 36482 39172 36484
rect 39116 36430 39118 36482
rect 39118 36430 39170 36482
rect 39170 36430 39172 36482
rect 39116 36428 39172 36430
rect 40348 46620 40404 46676
rect 40012 45276 40068 45332
rect 41580 46786 41636 46788
rect 41580 46734 41582 46786
rect 41582 46734 41634 46786
rect 41634 46734 41636 46786
rect 41580 46732 41636 46734
rect 41244 46674 41300 46676
rect 41244 46622 41246 46674
rect 41246 46622 41298 46674
rect 41298 46622 41300 46674
rect 41244 46620 41300 46622
rect 39788 44044 39844 44100
rect 40684 44268 40740 44324
rect 41132 44268 41188 44324
rect 40012 43708 40068 43764
rect 40348 44098 40404 44100
rect 40348 44046 40350 44098
rect 40350 44046 40402 44098
rect 40402 44046 40404 44098
rect 40348 44044 40404 44046
rect 39788 43426 39844 43428
rect 39788 43374 39790 43426
rect 39790 43374 39842 43426
rect 39842 43374 39844 43426
rect 39788 43372 39844 43374
rect 41132 42924 41188 42980
rect 40348 42700 40404 42756
rect 40124 41244 40180 41300
rect 39676 40572 39732 40628
rect 40124 40572 40180 40628
rect 42700 50540 42756 50596
rect 42364 50482 42420 50484
rect 42364 50430 42366 50482
rect 42366 50430 42418 50482
rect 42418 50430 42420 50482
rect 42364 50428 42420 50430
rect 42028 49868 42084 49924
rect 42364 49868 42420 49924
rect 43036 50594 43092 50596
rect 43036 50542 43038 50594
rect 43038 50542 43090 50594
rect 43090 50542 43092 50594
rect 43036 50540 43092 50542
rect 43372 50540 43428 50596
rect 42252 48914 42308 48916
rect 42252 48862 42254 48914
rect 42254 48862 42306 48914
rect 42306 48862 42308 48914
rect 42252 48860 42308 48862
rect 42028 48748 42084 48804
rect 42476 48802 42532 48804
rect 42476 48750 42478 48802
rect 42478 48750 42530 48802
rect 42530 48750 42532 48802
rect 42476 48748 42532 48750
rect 42700 48860 42756 48916
rect 42364 47628 42420 47684
rect 41804 46956 41860 47012
rect 42588 47458 42644 47460
rect 42588 47406 42590 47458
rect 42590 47406 42642 47458
rect 42642 47406 42644 47458
rect 42588 47404 42644 47406
rect 43148 47628 43204 47684
rect 42812 47234 42868 47236
rect 42812 47182 42814 47234
rect 42814 47182 42866 47234
rect 42866 47182 42868 47234
rect 42812 47180 42868 47182
rect 41804 46732 41860 46788
rect 41804 46396 41860 46452
rect 42588 46732 42644 46788
rect 42924 46620 42980 46676
rect 43036 46562 43092 46564
rect 43036 46510 43038 46562
rect 43038 46510 43090 46562
rect 43090 46510 43092 46562
rect 43036 46508 43092 46510
rect 42812 45890 42868 45892
rect 42812 45838 42814 45890
rect 42814 45838 42866 45890
rect 42866 45838 42868 45890
rect 42812 45836 42868 45838
rect 45724 50594 45780 50596
rect 45724 50542 45726 50594
rect 45726 50542 45778 50594
rect 45778 50542 45780 50594
rect 45724 50540 45780 50542
rect 43484 49922 43540 49924
rect 43484 49870 43486 49922
rect 43486 49870 43538 49922
rect 43538 49870 43540 49922
rect 43484 49868 43540 49870
rect 46060 49756 46116 49812
rect 45500 47404 45556 47460
rect 43372 46674 43428 46676
rect 43372 46622 43374 46674
rect 43374 46622 43426 46674
rect 43426 46622 43428 46674
rect 43372 46620 43428 46622
rect 45276 46620 45332 46676
rect 44156 46562 44212 46564
rect 44156 46510 44158 46562
rect 44158 46510 44210 46562
rect 44210 46510 44212 46562
rect 44156 46508 44212 46510
rect 42364 45164 42420 45220
rect 41916 45052 41972 45108
rect 41356 43596 41412 43652
rect 41468 43538 41524 43540
rect 41468 43486 41470 43538
rect 41470 43486 41522 43538
rect 41522 43486 41524 43538
rect 41468 43484 41524 43486
rect 41468 42924 41524 42980
rect 41020 41970 41076 41972
rect 41020 41918 41022 41970
rect 41022 41918 41074 41970
rect 41074 41918 41076 41970
rect 41020 41916 41076 41918
rect 40908 40626 40964 40628
rect 40908 40574 40910 40626
rect 40910 40574 40962 40626
rect 40962 40574 40964 40626
rect 40908 40572 40964 40574
rect 41244 40236 41300 40292
rect 38332 36258 38388 36260
rect 38332 36206 38334 36258
rect 38334 36206 38386 36258
rect 38386 36206 38388 36258
rect 38332 36204 38388 36206
rect 38220 35586 38276 35588
rect 38220 35534 38222 35586
rect 38222 35534 38274 35586
rect 38274 35534 38276 35586
rect 38220 35532 38276 35534
rect 37884 35084 37940 35140
rect 37436 34972 37492 35028
rect 38892 36258 38948 36260
rect 38892 36206 38894 36258
rect 38894 36206 38946 36258
rect 38946 36206 38948 36258
rect 38892 36204 38948 36206
rect 38892 35698 38948 35700
rect 38892 35646 38894 35698
rect 38894 35646 38946 35698
rect 38946 35646 38948 35698
rect 38892 35644 38948 35646
rect 38780 35196 38836 35252
rect 39004 35084 39060 35140
rect 39452 35644 39508 35700
rect 38780 34972 38836 35028
rect 38444 34524 38500 34580
rect 38556 34636 38612 34692
rect 37884 34354 37940 34356
rect 37884 34302 37886 34354
rect 37886 34302 37938 34354
rect 37938 34302 37940 34354
rect 37884 34300 37940 34302
rect 39228 34972 39284 35028
rect 38780 34636 38836 34692
rect 38780 34300 38836 34356
rect 38668 34242 38724 34244
rect 38668 34190 38670 34242
rect 38670 34190 38722 34242
rect 38722 34190 38724 34242
rect 38668 34188 38724 34190
rect 37548 33628 37604 33684
rect 37436 33404 37492 33460
rect 37772 32620 37828 32676
rect 37884 32396 37940 32452
rect 37100 29372 37156 29428
rect 36540 28642 36596 28644
rect 36540 28590 36542 28642
rect 36542 28590 36594 28642
rect 36594 28590 36596 28642
rect 36540 28588 36596 28590
rect 37324 28700 37380 28756
rect 37212 28642 37268 28644
rect 37212 28590 37214 28642
rect 37214 28590 37266 28642
rect 37266 28590 37268 28642
rect 37212 28588 37268 28590
rect 38556 34130 38612 34132
rect 38556 34078 38558 34130
rect 38558 34078 38610 34130
rect 38610 34078 38612 34130
rect 38556 34076 38612 34078
rect 38444 33628 38500 33684
rect 38108 33068 38164 33124
rect 37996 28588 38052 28644
rect 35980 27468 36036 27524
rect 35868 27020 35924 27076
rect 34860 26962 34916 26964
rect 34860 26910 34862 26962
rect 34862 26910 34914 26962
rect 34914 26910 34916 26962
rect 34860 26908 34916 26910
rect 36092 27132 36148 27188
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34860 25730 34916 25732
rect 34860 25678 34862 25730
rect 34862 25678 34914 25730
rect 34914 25678 34916 25730
rect 34860 25676 34916 25678
rect 34748 25282 34804 25284
rect 34748 25230 34750 25282
rect 34750 25230 34802 25282
rect 34802 25230 34804 25282
rect 34748 25228 34804 25230
rect 35084 25564 35140 25620
rect 34972 25116 35028 25172
rect 34412 23884 34468 23940
rect 34636 24610 34692 24612
rect 34636 24558 34638 24610
rect 34638 24558 34690 24610
rect 34690 24558 34692 24610
rect 34636 24556 34692 24558
rect 34972 23996 35028 24052
rect 34300 21308 34356 21364
rect 34300 20076 34356 20132
rect 34748 21756 34804 21812
rect 34860 21586 34916 21588
rect 34860 21534 34862 21586
rect 34862 21534 34914 21586
rect 34914 21534 34916 21586
rect 34860 21532 34916 21534
rect 35532 25228 35588 25284
rect 35532 24722 35588 24724
rect 35532 24670 35534 24722
rect 35534 24670 35586 24722
rect 35586 24670 35588 24722
rect 35532 24668 35588 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35308 21698 35364 21700
rect 35308 21646 35310 21698
rect 35310 21646 35362 21698
rect 35362 21646 35364 21698
rect 35308 21644 35364 21646
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34748 19964 34804 20020
rect 34524 19180 34580 19236
rect 34300 18844 34356 18900
rect 34076 18620 34132 18676
rect 32732 17164 32788 17220
rect 34188 17442 34244 17444
rect 34188 17390 34190 17442
rect 34190 17390 34242 17442
rect 34242 17390 34244 17442
rect 34188 17388 34244 17390
rect 33180 17276 33236 17332
rect 32060 15260 32116 15316
rect 31052 14812 31108 14868
rect 31164 14924 31220 14980
rect 31500 14306 31556 14308
rect 31500 14254 31502 14306
rect 31502 14254 31554 14306
rect 31554 14254 31556 14306
rect 31500 14252 31556 14254
rect 32508 15202 32564 15204
rect 32508 15150 32510 15202
rect 32510 15150 32562 15202
rect 32562 15150 32564 15202
rect 32508 15148 32564 15150
rect 31836 13020 31892 13076
rect 34188 16828 34244 16884
rect 33404 15148 33460 15204
rect 33740 15148 33796 15204
rect 33180 13132 33236 13188
rect 33628 12908 33684 12964
rect 33852 12124 33908 12180
rect 30828 10780 30884 10836
rect 31612 11394 31668 11396
rect 31612 11342 31614 11394
rect 31614 11342 31666 11394
rect 31666 11342 31668 11394
rect 31612 11340 31668 11342
rect 31948 11340 32004 11396
rect 31164 10668 31220 10724
rect 32620 11394 32676 11396
rect 32620 11342 32622 11394
rect 32622 11342 32674 11394
rect 32674 11342 32676 11394
rect 32620 11340 32676 11342
rect 32844 11228 32900 11284
rect 32396 11170 32452 11172
rect 32396 11118 32398 11170
rect 32398 11118 32450 11170
rect 32450 11118 32452 11170
rect 32396 11116 32452 11118
rect 33404 11116 33460 11172
rect 29036 8316 29092 8372
rect 28700 7980 28756 8036
rect 29484 7308 29540 7364
rect 31164 7698 31220 7700
rect 31164 7646 31166 7698
rect 31166 7646 31218 7698
rect 31218 7646 31220 7698
rect 31164 7644 31220 7646
rect 30828 7308 30884 7364
rect 30940 7250 30996 7252
rect 30940 7198 30942 7250
rect 30942 7198 30994 7250
rect 30994 7198 30996 7250
rect 30940 7196 30996 7198
rect 31052 6972 31108 7028
rect 31164 7308 31220 7364
rect 27804 6412 27860 6468
rect 27468 6130 27524 6132
rect 27468 6078 27470 6130
rect 27470 6078 27522 6130
rect 27522 6078 27524 6130
rect 27468 6076 27524 6078
rect 30380 6466 30436 6468
rect 30380 6414 30382 6466
rect 30382 6414 30434 6466
rect 30434 6414 30436 6466
rect 30380 6412 30436 6414
rect 31052 6466 31108 6468
rect 31052 6414 31054 6466
rect 31054 6414 31106 6466
rect 31106 6414 31108 6466
rect 31052 6412 31108 6414
rect 27692 5906 27748 5908
rect 27692 5854 27694 5906
rect 27694 5854 27746 5906
rect 27746 5854 27748 5906
rect 27692 5852 27748 5854
rect 27804 5122 27860 5124
rect 27804 5070 27806 5122
rect 27806 5070 27858 5122
rect 27858 5070 27860 5122
rect 27804 5068 27860 5070
rect 28476 5122 28532 5124
rect 28476 5070 28478 5122
rect 28478 5070 28530 5122
rect 28530 5070 28532 5122
rect 28476 5068 28532 5070
rect 28252 4898 28308 4900
rect 28252 4846 28254 4898
rect 28254 4846 28306 4898
rect 28306 4846 28308 4898
rect 28252 4844 28308 4846
rect 29932 4844 29988 4900
rect 33404 10332 33460 10388
rect 32172 9660 32228 9716
rect 31948 9154 32004 9156
rect 31948 9102 31950 9154
rect 31950 9102 32002 9154
rect 32002 9102 32004 9154
rect 31948 9100 32004 9102
rect 33068 9100 33124 9156
rect 33516 10444 33572 10500
rect 31724 8818 31780 8820
rect 31724 8766 31726 8818
rect 31726 8766 31778 8818
rect 31778 8766 31780 8818
rect 31724 8764 31780 8766
rect 33068 8818 33124 8820
rect 33068 8766 33070 8818
rect 33070 8766 33122 8818
rect 33122 8766 33124 8818
rect 33068 8764 33124 8766
rect 31388 8092 31444 8148
rect 31836 7698 31892 7700
rect 31836 7646 31838 7698
rect 31838 7646 31890 7698
rect 31890 7646 31892 7698
rect 31836 7644 31892 7646
rect 31388 6860 31444 6916
rect 32844 6914 32900 6916
rect 32844 6862 32846 6914
rect 32846 6862 32898 6914
rect 32898 6862 32900 6914
rect 32844 6860 32900 6862
rect 33628 9100 33684 9156
rect 34300 15820 34356 15876
rect 34748 12908 34804 12964
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35644 23938 35700 23940
rect 35644 23886 35646 23938
rect 35646 23886 35698 23938
rect 35698 23886 35700 23938
rect 35644 23884 35700 23886
rect 35980 23826 36036 23828
rect 35980 23774 35982 23826
rect 35982 23774 36034 23826
rect 36034 23774 36036 23826
rect 35980 23772 36036 23774
rect 36316 27074 36372 27076
rect 36316 27022 36318 27074
rect 36318 27022 36370 27074
rect 36370 27022 36372 27074
rect 36316 27020 36372 27022
rect 36428 25564 36484 25620
rect 36316 25116 36372 25172
rect 37100 27298 37156 27300
rect 37100 27246 37102 27298
rect 37102 27246 37154 27298
rect 37154 27246 37156 27298
rect 37100 27244 37156 27246
rect 37212 27074 37268 27076
rect 37212 27022 37214 27074
rect 37214 27022 37266 27074
rect 37266 27022 37268 27074
rect 37212 27020 37268 27022
rect 37660 26962 37716 26964
rect 37660 26910 37662 26962
rect 37662 26910 37714 26962
rect 37714 26910 37716 26962
rect 37660 26908 37716 26910
rect 37100 26850 37156 26852
rect 37100 26798 37102 26850
rect 37102 26798 37154 26850
rect 37154 26798 37156 26850
rect 37100 26796 37156 26798
rect 38108 27692 38164 27748
rect 37884 26850 37940 26852
rect 37884 26798 37886 26850
rect 37886 26798 37938 26850
rect 37938 26798 37940 26850
rect 37884 26796 37940 26798
rect 37212 23938 37268 23940
rect 37212 23886 37214 23938
rect 37214 23886 37266 23938
rect 37266 23886 37268 23938
rect 37212 23884 37268 23886
rect 36876 23826 36932 23828
rect 36876 23774 36878 23826
rect 36878 23774 36930 23826
rect 36930 23774 36932 23826
rect 36876 23772 36932 23774
rect 36764 23100 36820 23156
rect 37100 23714 37156 23716
rect 37100 23662 37102 23714
rect 37102 23662 37154 23714
rect 37154 23662 37156 23714
rect 37100 23660 37156 23662
rect 35644 21644 35700 21700
rect 35644 21420 35700 21476
rect 36092 21532 36148 21588
rect 35420 17724 35476 17780
rect 35980 20636 36036 20692
rect 35980 16716 36036 16772
rect 36204 21474 36260 21476
rect 36204 21422 36206 21474
rect 36206 21422 36258 21474
rect 36258 21422 36260 21474
rect 36204 21420 36260 21422
rect 36428 18956 36484 19012
rect 37996 24780 38052 24836
rect 37996 24556 38052 24612
rect 37212 22930 37268 22932
rect 37212 22878 37214 22930
rect 37214 22878 37266 22930
rect 37266 22878 37268 22930
rect 37212 22876 37268 22878
rect 37100 22428 37156 22484
rect 37100 21308 37156 21364
rect 37772 21586 37828 21588
rect 37772 21534 37774 21586
rect 37774 21534 37826 21586
rect 37826 21534 37828 21586
rect 37772 21532 37828 21534
rect 37772 20860 37828 20916
rect 37660 20748 37716 20804
rect 37324 20690 37380 20692
rect 37324 20638 37326 20690
rect 37326 20638 37378 20690
rect 37378 20638 37380 20690
rect 37324 20636 37380 20638
rect 38108 23436 38164 23492
rect 37100 19852 37156 19908
rect 37772 19404 37828 19460
rect 38668 32786 38724 32788
rect 38668 32734 38670 32786
rect 38670 32734 38722 32786
rect 38722 32734 38724 32786
rect 38668 32732 38724 32734
rect 39116 34860 39172 34916
rect 39004 34690 39060 34692
rect 39004 34638 39006 34690
rect 39006 34638 39058 34690
rect 39058 34638 39060 34690
rect 39004 34636 39060 34638
rect 41356 38834 41412 38836
rect 41356 38782 41358 38834
rect 41358 38782 41410 38834
rect 41410 38782 41412 38834
rect 41356 38780 41412 38782
rect 40236 36876 40292 36932
rect 40572 36482 40628 36484
rect 40572 36430 40574 36482
rect 40574 36430 40626 36482
rect 40626 36430 40628 36482
rect 40572 36428 40628 36430
rect 40236 35868 40292 35924
rect 40124 35308 40180 35364
rect 39788 34914 39844 34916
rect 39788 34862 39790 34914
rect 39790 34862 39842 34914
rect 39842 34862 39844 34914
rect 39788 34860 39844 34862
rect 39228 32844 39284 32900
rect 39116 32786 39172 32788
rect 39116 32734 39118 32786
rect 39118 32734 39170 32786
rect 39170 32734 39172 32786
rect 39116 32732 39172 32734
rect 39340 32396 39396 32452
rect 38780 28588 38836 28644
rect 39228 31948 39284 32004
rect 39004 30828 39060 30884
rect 39228 31724 39284 31780
rect 39564 34412 39620 34468
rect 40012 34860 40068 34916
rect 40236 34860 40292 34916
rect 41244 35756 41300 35812
rect 40236 34690 40292 34692
rect 40236 34638 40238 34690
rect 40238 34638 40290 34690
rect 40290 34638 40292 34690
rect 40236 34636 40292 34638
rect 40012 34412 40068 34468
rect 40124 31948 40180 32004
rect 39900 31778 39956 31780
rect 39900 31726 39902 31778
rect 39902 31726 39954 31778
rect 39954 31726 39956 31778
rect 39900 31724 39956 31726
rect 39564 31500 39620 31556
rect 41580 34748 41636 34804
rect 41244 33068 41300 33124
rect 41580 33964 41636 34020
rect 41692 33346 41748 33348
rect 41692 33294 41694 33346
rect 41694 33294 41746 33346
rect 41746 33294 41748 33346
rect 41692 33292 41748 33294
rect 41580 32956 41636 33012
rect 42476 45052 42532 45108
rect 43820 45276 43876 45332
rect 44268 45276 44324 45332
rect 44156 45164 44212 45220
rect 43708 44940 43764 44996
rect 45052 44322 45108 44324
rect 45052 44270 45054 44322
rect 45054 44270 45106 44322
rect 45106 44270 45108 44322
rect 45052 44268 45108 44270
rect 44268 44156 44324 44212
rect 44940 44210 44996 44212
rect 44940 44158 44942 44210
rect 44942 44158 44994 44210
rect 44994 44158 44996 44210
rect 44940 44156 44996 44158
rect 43708 43708 43764 43764
rect 42588 43484 42644 43540
rect 43484 43596 43540 43652
rect 41916 42252 41972 42308
rect 42588 41244 42644 41300
rect 41916 40514 41972 40516
rect 41916 40462 41918 40514
rect 41918 40462 41970 40514
rect 41970 40462 41972 40514
rect 41916 40460 41972 40462
rect 42028 40402 42084 40404
rect 42028 40350 42030 40402
rect 42030 40350 42082 40402
rect 42082 40350 42084 40402
rect 42028 40348 42084 40350
rect 43484 41298 43540 41300
rect 43484 41246 43486 41298
rect 43486 41246 43538 41298
rect 43538 41246 43540 41298
rect 43484 41244 43540 41246
rect 43036 40460 43092 40516
rect 43148 40908 43204 40964
rect 43036 36428 43092 36484
rect 42924 35756 42980 35812
rect 42140 35698 42196 35700
rect 42140 35646 42142 35698
rect 42142 35646 42194 35698
rect 42194 35646 42196 35698
rect 42140 35644 42196 35646
rect 42252 34748 42308 34804
rect 42812 35420 42868 35476
rect 44492 43650 44548 43652
rect 44492 43598 44494 43650
rect 44494 43598 44546 43650
rect 44546 43598 44548 43650
rect 44492 43596 44548 43598
rect 43932 40460 43988 40516
rect 43708 39004 43764 39060
rect 43820 38780 43876 38836
rect 43708 36482 43764 36484
rect 43708 36430 43710 36482
rect 43710 36430 43762 36482
rect 43762 36430 43764 36482
rect 43708 36428 43764 36430
rect 44156 40962 44212 40964
rect 44156 40910 44158 40962
rect 44158 40910 44210 40962
rect 44210 40910 44212 40962
rect 44156 40908 44212 40910
rect 44044 40348 44100 40404
rect 44940 42028 44996 42084
rect 45052 41804 45108 41860
rect 49196 50540 49252 50596
rect 48972 49922 49028 49924
rect 48972 49870 48974 49922
rect 48974 49870 49026 49922
rect 49026 49870 49028 49922
rect 48972 49868 49028 49870
rect 48860 49810 48916 49812
rect 48860 49758 48862 49810
rect 48862 49758 48914 49810
rect 48914 49758 48916 49810
rect 48860 49756 48916 49758
rect 49756 50540 49812 50596
rect 49980 50428 50036 50484
rect 51212 50428 51268 50484
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 46620 48802 46676 48804
rect 46620 48750 46622 48802
rect 46622 48750 46674 48802
rect 46674 48750 46676 48802
rect 46620 48748 46676 48750
rect 47180 48748 47236 48804
rect 47180 48354 47236 48356
rect 47180 48302 47182 48354
rect 47182 48302 47234 48354
rect 47234 48302 47236 48354
rect 47180 48300 47236 48302
rect 46508 48076 46564 48132
rect 46620 47964 46676 48020
rect 47404 48076 47460 48132
rect 48188 48130 48244 48132
rect 48188 48078 48190 48130
rect 48190 48078 48242 48130
rect 48242 48078 48244 48130
rect 48188 48076 48244 48078
rect 45948 47068 46004 47124
rect 47740 48018 47796 48020
rect 47740 47966 47742 48018
rect 47742 47966 47794 48018
rect 47794 47966 47796 48018
rect 47740 47964 47796 47966
rect 47740 47404 47796 47460
rect 45836 46284 45892 46340
rect 46284 45612 46340 45668
rect 45612 44322 45668 44324
rect 45612 44270 45614 44322
rect 45614 44270 45666 44322
rect 45666 44270 45668 44322
rect 45612 44268 45668 44270
rect 46620 45276 46676 45332
rect 47740 46284 47796 46340
rect 47068 44828 47124 44884
rect 45388 43596 45444 43652
rect 46060 43596 46116 43652
rect 45164 40290 45220 40292
rect 45164 40238 45166 40290
rect 45166 40238 45218 40290
rect 45218 40238 45220 40290
rect 45164 40236 45220 40238
rect 44044 39452 44100 39508
rect 44380 39058 44436 39060
rect 44380 39006 44382 39058
rect 44382 39006 44434 39058
rect 44434 39006 44436 39058
rect 44380 39004 44436 39006
rect 44828 39506 44884 39508
rect 44828 39454 44830 39506
rect 44830 39454 44882 39506
rect 44882 39454 44884 39506
rect 44828 39452 44884 39454
rect 44940 39116 44996 39172
rect 44044 38668 44100 38724
rect 44380 37660 44436 37716
rect 43596 35420 43652 35476
rect 43708 35308 43764 35364
rect 43932 35308 43988 35364
rect 43372 35196 43428 35252
rect 42476 34802 42532 34804
rect 42476 34750 42478 34802
rect 42478 34750 42530 34802
rect 42530 34750 42532 34802
rect 42476 34748 42532 34750
rect 42028 33292 42084 33348
rect 42140 33068 42196 33124
rect 40348 31164 40404 31220
rect 39452 29986 39508 29988
rect 39452 29934 39454 29986
rect 39454 29934 39506 29986
rect 39506 29934 39508 29986
rect 39452 29932 39508 29934
rect 39340 29708 39396 29764
rect 39228 29650 39284 29652
rect 39228 29598 39230 29650
rect 39230 29598 39282 29650
rect 39282 29598 39284 29650
rect 39228 29596 39284 29598
rect 39004 28588 39060 28644
rect 39004 28252 39060 28308
rect 39116 28028 39172 28084
rect 38556 27692 38612 27748
rect 38444 26908 38500 26964
rect 38332 26066 38388 26068
rect 38332 26014 38334 26066
rect 38334 26014 38386 26066
rect 38386 26014 38388 26066
rect 38332 26012 38388 26014
rect 38332 25564 38388 25620
rect 38332 23660 38388 23716
rect 39116 26908 39172 26964
rect 40572 29986 40628 29988
rect 40572 29934 40574 29986
rect 40574 29934 40626 29986
rect 40626 29934 40628 29986
rect 40572 29932 40628 29934
rect 39900 29314 39956 29316
rect 39900 29262 39902 29314
rect 39902 29262 39954 29314
rect 39954 29262 39956 29314
rect 39900 29260 39956 29262
rect 40012 29036 40068 29092
rect 39452 28252 39508 28308
rect 39340 27692 39396 27748
rect 39564 28028 39620 28084
rect 39228 27020 39284 27076
rect 38780 24668 38836 24724
rect 39004 24722 39060 24724
rect 39004 24670 39006 24722
rect 39006 24670 39058 24722
rect 39058 24670 39060 24722
rect 39004 24668 39060 24670
rect 38556 23884 38612 23940
rect 38668 21756 38724 21812
rect 36540 17778 36596 17780
rect 36540 17726 36542 17778
rect 36542 17726 36594 17778
rect 36594 17726 36596 17778
rect 36540 17724 36596 17726
rect 36428 17388 36484 17444
rect 36652 17164 36708 17220
rect 36316 16716 36372 16772
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35308 15538 35364 15540
rect 35308 15486 35310 15538
rect 35310 15486 35362 15538
rect 35362 15486 35364 15538
rect 35308 15484 35364 15486
rect 36204 15820 36260 15876
rect 35644 15260 35700 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35980 13804 36036 13860
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13020 35700 13076
rect 34860 12572 34916 12628
rect 35644 12684 35700 12740
rect 34748 12178 34804 12180
rect 34748 12126 34750 12178
rect 34750 12126 34802 12178
rect 34802 12126 34804 12178
rect 34748 12124 34804 12126
rect 35980 12348 36036 12404
rect 36092 12796 36148 12852
rect 36204 12684 36260 12740
rect 36428 15484 36484 15540
rect 36652 13746 36708 13748
rect 36652 13694 36654 13746
rect 36654 13694 36706 13746
rect 36706 13694 36708 13746
rect 36652 13692 36708 13694
rect 36428 12738 36484 12740
rect 36428 12686 36430 12738
rect 36430 12686 36482 12738
rect 36482 12686 36484 12738
rect 36428 12684 36484 12686
rect 36316 12290 36372 12292
rect 36316 12238 36318 12290
rect 36318 12238 36370 12290
rect 36370 12238 36372 12290
rect 36316 12236 36372 12238
rect 34300 11340 34356 11396
rect 35196 12012 35252 12068
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35084 11228 35140 11284
rect 35644 10892 35700 10948
rect 35868 10780 35924 10836
rect 35756 10668 35812 10724
rect 35644 10332 35700 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35532 9548 35588 9604
rect 35644 9266 35700 9268
rect 35644 9214 35646 9266
rect 35646 9214 35698 9266
rect 35698 9214 35700 9266
rect 35644 9212 35700 9214
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35420 8316 35476 8372
rect 34972 8146 35028 8148
rect 34972 8094 34974 8146
rect 34974 8094 35026 8146
rect 35026 8094 35028 8146
rect 34972 8092 35028 8094
rect 36428 11564 36484 11620
rect 36204 10668 36260 10724
rect 35980 10498 36036 10500
rect 35980 10446 35982 10498
rect 35982 10446 36034 10498
rect 36034 10446 36036 10498
rect 35980 10444 36036 10446
rect 36204 10108 36260 10164
rect 35980 9548 36036 9604
rect 35868 9154 35924 9156
rect 35868 9102 35870 9154
rect 35870 9102 35922 9154
rect 35922 9102 35924 9154
rect 35868 9100 35924 9102
rect 36764 10722 36820 10724
rect 36764 10670 36766 10722
rect 36766 10670 36818 10722
rect 36818 10670 36820 10722
rect 36764 10668 36820 10670
rect 36428 9266 36484 9268
rect 36428 9214 36430 9266
rect 36430 9214 36482 9266
rect 36482 9214 36484 9266
rect 36428 9212 36484 9214
rect 36876 9212 36932 9268
rect 35756 8316 35812 8372
rect 35644 8258 35700 8260
rect 35644 8206 35646 8258
rect 35646 8206 35698 8258
rect 35698 8206 35700 8258
rect 35644 8204 35700 8206
rect 36316 8370 36372 8372
rect 36316 8318 36318 8370
rect 36318 8318 36370 8370
rect 36370 8318 36372 8370
rect 36316 8316 36372 8318
rect 35756 8146 35812 8148
rect 35756 8094 35758 8146
rect 35758 8094 35810 8146
rect 35810 8094 35812 8146
rect 35756 8092 35812 8094
rect 36540 8092 36596 8148
rect 34188 7644 34244 7700
rect 31276 5068 31332 5124
rect 33404 5180 33460 5236
rect 36092 7586 36148 7588
rect 36092 7534 36094 7586
rect 36094 7534 36146 7586
rect 36146 7534 36148 7586
rect 36092 7532 36148 7534
rect 39340 27356 39396 27412
rect 39340 24610 39396 24612
rect 39340 24558 39342 24610
rect 39342 24558 39394 24610
rect 39394 24558 39396 24610
rect 39340 24556 39396 24558
rect 40460 29372 40516 29428
rect 40012 28028 40068 28084
rect 40236 28418 40292 28420
rect 40236 28366 40238 28418
rect 40238 28366 40290 28418
rect 40290 28366 40292 28418
rect 40236 28364 40292 28366
rect 40236 28082 40292 28084
rect 40236 28030 40238 28082
rect 40238 28030 40290 28082
rect 40290 28030 40292 28082
rect 40236 28028 40292 28030
rect 41132 29426 41188 29428
rect 41132 29374 41134 29426
rect 41134 29374 41186 29426
rect 41186 29374 41188 29426
rect 41132 29372 41188 29374
rect 40572 28588 40628 28644
rect 39676 27356 39732 27412
rect 40236 27468 40292 27524
rect 40012 26962 40068 26964
rect 40012 26910 40014 26962
rect 40014 26910 40066 26962
rect 40066 26910 40068 26962
rect 40012 26908 40068 26910
rect 40348 26908 40404 26964
rect 39900 26460 39956 26516
rect 40012 26572 40068 26628
rect 39900 26178 39956 26180
rect 39900 26126 39902 26178
rect 39902 26126 39954 26178
rect 39954 26126 39956 26178
rect 39900 26124 39956 26126
rect 39676 25116 39732 25172
rect 39788 23436 39844 23492
rect 39452 23266 39508 23268
rect 39452 23214 39454 23266
rect 39454 23214 39506 23266
rect 39506 23214 39508 23266
rect 39452 23212 39508 23214
rect 39116 22876 39172 22932
rect 39676 22930 39732 22932
rect 39676 22878 39678 22930
rect 39678 22878 39730 22930
rect 39730 22878 39732 22930
rect 39676 22876 39732 22878
rect 39788 21756 39844 21812
rect 39116 20802 39172 20804
rect 39116 20750 39118 20802
rect 39118 20750 39170 20802
rect 39170 20750 39172 20802
rect 39116 20748 39172 20750
rect 39900 20188 39956 20244
rect 40012 23548 40068 23604
rect 39228 20076 39284 20132
rect 37324 15314 37380 15316
rect 37324 15262 37326 15314
rect 37326 15262 37378 15314
rect 37378 15262 37380 15314
rect 37324 15260 37380 15262
rect 38220 17500 38276 17556
rect 37548 17388 37604 17444
rect 37996 17106 38052 17108
rect 37996 17054 37998 17106
rect 37998 17054 38050 17106
rect 38050 17054 38052 17106
rect 37996 17052 38052 17054
rect 38108 16828 38164 16884
rect 37660 15874 37716 15876
rect 37660 15822 37662 15874
rect 37662 15822 37714 15874
rect 37714 15822 37716 15874
rect 37660 15820 37716 15822
rect 38220 14476 38276 14532
rect 37548 13132 37604 13188
rect 37436 12908 37492 12964
rect 37324 11676 37380 11732
rect 37324 10834 37380 10836
rect 37324 10782 37326 10834
rect 37326 10782 37378 10834
rect 37378 10782 37380 10834
rect 37324 10780 37380 10782
rect 38332 16492 38388 16548
rect 38556 17442 38612 17444
rect 38556 17390 38558 17442
rect 38558 17390 38610 17442
rect 38610 17390 38612 17442
rect 38556 17388 38612 17390
rect 38780 19010 38836 19012
rect 38780 18958 38782 19010
rect 38782 18958 38834 19010
rect 38834 18958 38836 19010
rect 38780 18956 38836 18958
rect 39452 19964 39508 20020
rect 38892 17836 38948 17892
rect 38668 17164 38724 17220
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 38556 17052 38612 17108
rect 38668 16940 38724 16996
rect 38556 15708 38612 15764
rect 39004 16828 39060 16884
rect 39004 16098 39060 16100
rect 39004 16046 39006 16098
rect 39006 16046 39058 16098
rect 39058 16046 39060 16098
rect 39004 16044 39060 16046
rect 38780 15426 38836 15428
rect 38780 15374 38782 15426
rect 38782 15374 38834 15426
rect 38834 15374 38836 15426
rect 38780 15372 38836 15374
rect 38444 14364 38500 14420
rect 38332 12908 38388 12964
rect 37996 12236 38052 12292
rect 38108 12684 38164 12740
rect 38108 12178 38164 12180
rect 38108 12126 38110 12178
rect 38110 12126 38162 12178
rect 38162 12126 38164 12178
rect 38108 12124 38164 12126
rect 37884 11900 37940 11956
rect 39228 17554 39284 17556
rect 39228 17502 39230 17554
rect 39230 17502 39282 17554
rect 39282 17502 39284 17554
rect 39228 17500 39284 17502
rect 39788 20018 39844 20020
rect 39788 19966 39790 20018
rect 39790 19966 39842 20018
rect 39842 19966 39844 20018
rect 39788 19964 39844 19966
rect 40348 24722 40404 24724
rect 40348 24670 40350 24722
rect 40350 24670 40402 24722
rect 40402 24670 40404 24722
rect 40348 24668 40404 24670
rect 40684 27356 40740 27412
rect 40796 28476 40852 28532
rect 40684 27074 40740 27076
rect 40684 27022 40686 27074
rect 40686 27022 40738 27074
rect 40738 27022 40740 27074
rect 40684 27020 40740 27022
rect 41020 28364 41076 28420
rect 41020 28082 41076 28084
rect 41020 28030 41022 28082
rect 41022 28030 41074 28082
rect 41074 28030 41076 28082
rect 41020 28028 41076 28030
rect 40236 20748 40292 20804
rect 39564 19122 39620 19124
rect 39564 19070 39566 19122
rect 39566 19070 39618 19122
rect 39618 19070 39620 19122
rect 39564 19068 39620 19070
rect 39564 17388 39620 17444
rect 40572 21532 40628 21588
rect 41020 26962 41076 26964
rect 41020 26910 41022 26962
rect 41022 26910 41074 26962
rect 41074 26910 41076 26962
rect 41020 26908 41076 26910
rect 40796 25228 40852 25284
rect 41804 32562 41860 32564
rect 41804 32510 41806 32562
rect 41806 32510 41858 32562
rect 41858 32510 41860 32562
rect 41804 32508 41860 32510
rect 42588 34018 42644 34020
rect 42588 33966 42590 34018
rect 42590 33966 42642 34018
rect 42642 33966 42644 34018
rect 42588 33964 42644 33966
rect 42588 33628 42644 33684
rect 42476 33068 42532 33124
rect 42924 33964 42980 34020
rect 43036 33068 43092 33124
rect 44268 36204 44324 36260
rect 44268 35756 44324 35812
rect 43708 35084 43764 35140
rect 43484 33570 43540 33572
rect 43484 33518 43486 33570
rect 43486 33518 43538 33570
rect 43538 33518 43540 33570
rect 43484 33516 43540 33518
rect 43148 32844 43204 32900
rect 42028 32060 42084 32116
rect 43260 32508 43316 32564
rect 42140 31052 42196 31108
rect 42140 30268 42196 30324
rect 41356 29932 41412 29988
rect 42028 29596 42084 29652
rect 41356 28642 41412 28644
rect 41356 28590 41358 28642
rect 41358 28590 41410 28642
rect 41410 28590 41412 28642
rect 41356 28588 41412 28590
rect 41804 28530 41860 28532
rect 41804 28478 41806 28530
rect 41806 28478 41858 28530
rect 41858 28478 41860 28530
rect 41804 28476 41860 28478
rect 41468 27692 41524 27748
rect 41468 27074 41524 27076
rect 41468 27022 41470 27074
rect 41470 27022 41522 27074
rect 41522 27022 41524 27074
rect 41468 27020 41524 27022
rect 42812 31554 42868 31556
rect 42812 31502 42814 31554
rect 42814 31502 42866 31554
rect 42866 31502 42868 31554
rect 42812 31500 42868 31502
rect 42588 30156 42644 30212
rect 42700 29314 42756 29316
rect 42700 29262 42702 29314
rect 42702 29262 42754 29314
rect 42754 29262 42756 29314
rect 42700 29260 42756 29262
rect 42588 28812 42644 28868
rect 43148 30210 43204 30212
rect 43148 30158 43150 30210
rect 43150 30158 43202 30210
rect 43202 30158 43204 30210
rect 43148 30156 43204 30158
rect 42700 28476 42756 28532
rect 43148 29932 43204 29988
rect 41244 24892 41300 24948
rect 43036 26178 43092 26180
rect 43036 26126 43038 26178
rect 43038 26126 43090 26178
rect 43090 26126 43092 26178
rect 43036 26124 43092 26126
rect 40908 23548 40964 23604
rect 41244 24668 41300 24724
rect 41356 23212 41412 23268
rect 41244 22764 41300 22820
rect 41020 21362 41076 21364
rect 41020 21310 41022 21362
rect 41022 21310 41074 21362
rect 41074 21310 41076 21362
rect 41020 21308 41076 21310
rect 41020 21084 41076 21140
rect 41804 23212 41860 23268
rect 42700 23212 42756 23268
rect 42140 22988 42196 23044
rect 41804 22876 41860 22932
rect 41580 22146 41636 22148
rect 41580 22094 41582 22146
rect 41582 22094 41634 22146
rect 41634 22094 41636 22146
rect 41580 22092 41636 22094
rect 41580 21586 41636 21588
rect 41580 21534 41582 21586
rect 41582 21534 41634 21586
rect 41634 21534 41636 21586
rect 41580 21532 41636 21534
rect 42588 22876 42644 22932
rect 42476 21980 42532 22036
rect 42140 21756 42196 21812
rect 42364 21698 42420 21700
rect 42364 21646 42366 21698
rect 42366 21646 42418 21698
rect 42418 21646 42420 21698
rect 42364 21644 42420 21646
rect 41132 20076 41188 20132
rect 40348 18396 40404 18452
rect 40236 17164 40292 17220
rect 39452 16828 39508 16884
rect 39228 15932 39284 15988
rect 39340 16716 39396 16772
rect 39564 16492 39620 16548
rect 41244 19234 41300 19236
rect 41244 19182 41246 19234
rect 41246 19182 41298 19234
rect 41298 19182 41300 19234
rect 41244 19180 41300 19182
rect 41468 20860 41524 20916
rect 41580 20636 41636 20692
rect 41692 20578 41748 20580
rect 41692 20526 41694 20578
rect 41694 20526 41746 20578
rect 41746 20526 41748 20578
rect 41692 20524 41748 20526
rect 42028 20972 42084 21028
rect 41580 20076 41636 20132
rect 41468 20018 41524 20020
rect 41468 19966 41470 20018
rect 41470 19966 41522 20018
rect 41522 19966 41524 20018
rect 41468 19964 41524 19966
rect 41356 19068 41412 19124
rect 40908 18396 40964 18452
rect 40684 17778 40740 17780
rect 40684 17726 40686 17778
rect 40686 17726 40738 17778
rect 40738 17726 40740 17778
rect 40684 17724 40740 17726
rect 40572 17612 40628 17668
rect 40236 16940 40292 16996
rect 40236 16156 40292 16212
rect 40348 16268 40404 16324
rect 39788 15932 39844 15988
rect 39564 15820 39620 15876
rect 39004 13804 39060 13860
rect 38668 12402 38724 12404
rect 38668 12350 38670 12402
rect 38670 12350 38722 12402
rect 38722 12350 38724 12402
rect 38668 12348 38724 12350
rect 38780 12124 38836 12180
rect 38780 10668 38836 10724
rect 37772 10108 37828 10164
rect 38108 9154 38164 9156
rect 38108 9102 38110 9154
rect 38110 9102 38162 9154
rect 38162 9102 38164 9154
rect 38108 9100 38164 9102
rect 36988 8146 37044 8148
rect 36988 8094 36990 8146
rect 36990 8094 37042 8146
rect 37042 8094 37044 8146
rect 36988 8092 37044 8094
rect 36988 7474 37044 7476
rect 36988 7422 36990 7474
rect 36990 7422 37042 7474
rect 37042 7422 37044 7474
rect 36988 7420 37044 7422
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 37884 7586 37940 7588
rect 37884 7534 37886 7586
rect 37886 7534 37938 7586
rect 37938 7534 37940 7586
rect 37884 7532 37940 7534
rect 39116 13580 39172 13636
rect 40348 15708 40404 15764
rect 39676 14418 39732 14420
rect 39676 14366 39678 14418
rect 39678 14366 39730 14418
rect 39730 14366 39732 14418
rect 39676 14364 39732 14366
rect 40124 14364 40180 14420
rect 40124 13858 40180 13860
rect 40124 13806 40126 13858
rect 40126 13806 40178 13858
rect 40178 13806 40180 13858
rect 40124 13804 40180 13806
rect 39676 13746 39732 13748
rect 39676 13694 39678 13746
rect 39678 13694 39730 13746
rect 39730 13694 39732 13746
rect 39676 13692 39732 13694
rect 39116 12962 39172 12964
rect 39116 12910 39118 12962
rect 39118 12910 39170 12962
rect 39170 12910 39172 12962
rect 39116 12908 39172 12910
rect 39004 12012 39060 12068
rect 39004 11788 39060 11844
rect 38332 9266 38388 9268
rect 38332 9214 38334 9266
rect 38334 9214 38386 9266
rect 38386 9214 38388 9266
rect 38332 9212 38388 9214
rect 38668 9826 38724 9828
rect 38668 9774 38670 9826
rect 38670 9774 38722 9826
rect 38722 9774 38724 9826
rect 38668 9772 38724 9774
rect 37996 7474 38052 7476
rect 37996 7422 37998 7474
rect 37998 7422 38050 7474
rect 38050 7422 38052 7474
rect 37996 7420 38052 7422
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34076 5234 34132 5236
rect 34076 5182 34078 5234
rect 34078 5182 34130 5234
rect 34130 5182 34132 5234
rect 34076 5180 34132 5182
rect 33964 4956 34020 5012
rect 35420 4956 35476 5012
rect 37324 4956 37380 5012
rect 37996 4956 38052 5012
rect 38332 8540 38388 8596
rect 39116 10444 39172 10500
rect 39564 12850 39620 12852
rect 39564 12798 39566 12850
rect 39566 12798 39618 12850
rect 39618 12798 39620 12850
rect 39564 12796 39620 12798
rect 40124 12012 40180 12068
rect 40236 13356 40292 13412
rect 39900 11788 39956 11844
rect 39564 10722 39620 10724
rect 39564 10670 39566 10722
rect 39566 10670 39618 10722
rect 39618 10670 39620 10722
rect 39564 10668 39620 10670
rect 39452 10444 39508 10500
rect 39228 10050 39284 10052
rect 39228 9998 39230 10050
rect 39230 9998 39282 10050
rect 39282 9998 39284 10050
rect 39228 9996 39284 9998
rect 38892 8540 38948 8596
rect 39228 7868 39284 7924
rect 38780 7644 38836 7700
rect 38668 7586 38724 7588
rect 38668 7534 38670 7586
rect 38670 7534 38722 7586
rect 38722 7534 38724 7586
rect 38668 7532 38724 7534
rect 38332 6636 38388 6692
rect 39004 7698 39060 7700
rect 39004 7646 39006 7698
rect 39006 7646 39058 7698
rect 39058 7646 39060 7698
rect 39004 7644 39060 7646
rect 39676 10108 39732 10164
rect 39116 6690 39172 6692
rect 39116 6638 39118 6690
rect 39118 6638 39170 6690
rect 39170 6638 39172 6690
rect 39116 6636 39172 6638
rect 39228 5180 39284 5236
rect 38780 4338 38836 4340
rect 38780 4286 38782 4338
rect 38782 4286 38834 4338
rect 38834 4286 38836 4338
rect 38780 4284 38836 4286
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 30604 3500 30660 3556
rect 34076 3612 34132 3668
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 40460 12850 40516 12852
rect 40460 12798 40462 12850
rect 40462 12798 40514 12850
rect 40514 12798 40516 12850
rect 40460 12796 40516 12798
rect 40684 11788 40740 11844
rect 42140 20802 42196 20804
rect 42140 20750 42142 20802
rect 42142 20750 42194 20802
rect 42194 20750 42196 20802
rect 42140 20748 42196 20750
rect 42476 20188 42532 20244
rect 41804 20130 41860 20132
rect 41804 20078 41806 20130
rect 41806 20078 41858 20130
rect 41858 20078 41860 20130
rect 41804 20076 41860 20078
rect 41692 19180 41748 19236
rect 42140 19964 42196 20020
rect 41916 19068 41972 19124
rect 43372 31778 43428 31780
rect 43372 31726 43374 31778
rect 43374 31726 43426 31778
rect 43426 31726 43428 31778
rect 43372 31724 43428 31726
rect 44156 35532 44212 35588
rect 43372 31388 43428 31444
rect 43372 30268 43428 30324
rect 43932 32396 43988 32452
rect 43820 31836 43876 31892
rect 43820 31218 43876 31220
rect 43820 31166 43822 31218
rect 43822 31166 43874 31218
rect 43874 31166 43876 31218
rect 43820 31164 43876 31166
rect 43484 28812 43540 28868
rect 43708 27244 43764 27300
rect 43372 25282 43428 25284
rect 43372 25230 43374 25282
rect 43374 25230 43426 25282
rect 43426 25230 43428 25282
rect 43372 25228 43428 25230
rect 43820 29596 43876 29652
rect 43820 26124 43876 26180
rect 43708 25452 43764 25508
rect 44380 34690 44436 34692
rect 44380 34638 44382 34690
rect 44382 34638 44434 34690
rect 44434 34638 44436 34690
rect 44380 34636 44436 34638
rect 44380 34300 44436 34356
rect 44156 34130 44212 34132
rect 44156 34078 44158 34130
rect 44158 34078 44210 34130
rect 44210 34078 44212 34130
rect 44156 34076 44212 34078
rect 46732 43596 46788 43652
rect 47852 45276 47908 45332
rect 48972 48300 49028 48356
rect 49196 48130 49252 48132
rect 49196 48078 49198 48130
rect 49198 48078 49250 48130
rect 49250 48078 49252 48130
rect 49196 48076 49252 48078
rect 49084 47516 49140 47572
rect 51660 51378 51716 51380
rect 51660 51326 51662 51378
rect 51662 51326 51714 51378
rect 51714 51326 51716 51378
rect 51660 51324 51716 51326
rect 51436 50540 51492 50596
rect 49644 47570 49700 47572
rect 49644 47518 49646 47570
rect 49646 47518 49698 47570
rect 49698 47518 49700 47570
rect 49644 47516 49700 47518
rect 49532 47458 49588 47460
rect 49532 47406 49534 47458
rect 49534 47406 49586 47458
rect 49586 47406 49588 47458
rect 49532 47404 49588 47406
rect 48860 46508 48916 46564
rect 48748 46284 48804 46340
rect 48300 45948 48356 46004
rect 49196 45948 49252 46004
rect 49084 45500 49140 45556
rect 48748 45330 48804 45332
rect 48748 45278 48750 45330
rect 48750 45278 48802 45330
rect 48802 45278 48804 45330
rect 48748 45276 48804 45278
rect 47516 44828 47572 44884
rect 47068 42754 47124 42756
rect 47068 42702 47070 42754
rect 47070 42702 47122 42754
rect 47122 42702 47124 42754
rect 47068 42700 47124 42702
rect 46284 42028 46340 42084
rect 46732 41858 46788 41860
rect 46732 41806 46734 41858
rect 46734 41806 46786 41858
rect 46786 41806 46788 41858
rect 46732 41804 46788 41806
rect 51884 48860 51940 48916
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50428 46674 50484 46676
rect 50428 46622 50430 46674
rect 50430 46622 50482 46674
rect 50482 46622 50484 46674
rect 50428 46620 50484 46622
rect 48860 43260 48916 43316
rect 48524 43036 48580 43092
rect 47404 42700 47460 42756
rect 47964 41970 48020 41972
rect 47964 41918 47966 41970
rect 47966 41918 48018 41970
rect 48018 41918 48020 41970
rect 47964 41916 48020 41918
rect 49084 41970 49140 41972
rect 49084 41918 49086 41970
rect 49086 41918 49138 41970
rect 49138 41918 49140 41970
rect 49084 41916 49140 41918
rect 45500 38668 45556 38724
rect 46060 37884 46116 37940
rect 45164 37100 45220 37156
rect 44828 36482 44884 36484
rect 44828 36430 44830 36482
rect 44830 36430 44882 36482
rect 44882 36430 44884 36482
rect 44828 36428 44884 36430
rect 45836 37154 45892 37156
rect 45836 37102 45838 37154
rect 45838 37102 45890 37154
rect 45890 37102 45892 37154
rect 45836 37100 45892 37102
rect 45724 36594 45780 36596
rect 45724 36542 45726 36594
rect 45726 36542 45778 36594
rect 45778 36542 45780 36594
rect 45724 36540 45780 36542
rect 45164 36258 45220 36260
rect 45164 36206 45166 36258
rect 45166 36206 45218 36258
rect 45218 36206 45220 36258
rect 45164 36204 45220 36206
rect 44828 35810 44884 35812
rect 44828 35758 44830 35810
rect 44830 35758 44882 35810
rect 44882 35758 44884 35810
rect 44828 35756 44884 35758
rect 44156 32562 44212 32564
rect 44156 32510 44158 32562
rect 44158 32510 44210 32562
rect 44210 32510 44212 32562
rect 44156 32508 44212 32510
rect 45948 36370 46004 36372
rect 45948 36318 45950 36370
rect 45950 36318 46002 36370
rect 46002 36318 46004 36370
rect 45948 36316 46004 36318
rect 45276 35586 45332 35588
rect 45276 35534 45278 35586
rect 45278 35534 45330 35586
rect 45330 35534 45332 35586
rect 45276 35532 45332 35534
rect 45164 35026 45220 35028
rect 45164 34974 45166 35026
rect 45166 34974 45218 35026
rect 45218 34974 45220 35026
rect 45164 34972 45220 34974
rect 45276 34914 45332 34916
rect 45276 34862 45278 34914
rect 45278 34862 45330 34914
rect 45330 34862 45332 34914
rect 45276 34860 45332 34862
rect 46396 39116 46452 39172
rect 48524 40236 48580 40292
rect 49196 41074 49252 41076
rect 49196 41022 49198 41074
rect 49198 41022 49250 41074
rect 49250 41022 49252 41074
rect 49196 41020 49252 41022
rect 49196 39618 49252 39620
rect 49196 39566 49198 39618
rect 49198 39566 49250 39618
rect 49250 39566 49252 39618
rect 49196 39564 49252 39566
rect 46172 37100 46228 37156
rect 46732 35026 46788 35028
rect 46732 34974 46734 35026
rect 46734 34974 46786 35026
rect 46786 34974 46788 35026
rect 46732 34972 46788 34974
rect 45612 34802 45668 34804
rect 45612 34750 45614 34802
rect 45614 34750 45666 34802
rect 45666 34750 45668 34802
rect 45612 34748 45668 34750
rect 45052 34636 45108 34692
rect 45052 33740 45108 33796
rect 44492 33292 44548 33348
rect 45388 33346 45444 33348
rect 45388 33294 45390 33346
rect 45390 33294 45442 33346
rect 45442 33294 45444 33346
rect 45388 33292 45444 33294
rect 45052 33068 45108 33124
rect 45724 33122 45780 33124
rect 45724 33070 45726 33122
rect 45726 33070 45778 33122
rect 45778 33070 45780 33122
rect 45724 33068 45780 33070
rect 44940 32562 44996 32564
rect 44940 32510 44942 32562
rect 44942 32510 44994 32562
rect 44994 32510 44996 32562
rect 44940 32508 44996 32510
rect 44380 31052 44436 31108
rect 44828 31164 44884 31220
rect 45612 32562 45668 32564
rect 45612 32510 45614 32562
rect 45614 32510 45666 32562
rect 45666 32510 45668 32562
rect 45612 32508 45668 32510
rect 45052 32338 45108 32340
rect 45052 32286 45054 32338
rect 45054 32286 45106 32338
rect 45106 32286 45108 32338
rect 45052 32284 45108 32286
rect 46060 33346 46116 33348
rect 46060 33294 46062 33346
rect 46062 33294 46114 33346
rect 46114 33294 46116 33346
rect 46060 33292 46116 33294
rect 45276 31612 45332 31668
rect 45052 31106 45108 31108
rect 45052 31054 45054 31106
rect 45054 31054 45106 31106
rect 45106 31054 45108 31106
rect 45052 31052 45108 31054
rect 44268 27858 44324 27860
rect 44268 27806 44270 27858
rect 44270 27806 44322 27858
rect 44322 27806 44324 27858
rect 44268 27804 44324 27806
rect 44380 26796 44436 26852
rect 44268 26178 44324 26180
rect 44268 26126 44270 26178
rect 44270 26126 44322 26178
rect 44322 26126 44324 26178
rect 44268 26124 44324 26126
rect 44268 25452 44324 25508
rect 43820 24780 43876 24836
rect 43820 23548 43876 23604
rect 44044 24498 44100 24500
rect 44044 24446 44046 24498
rect 44046 24446 44098 24498
rect 44098 24446 44100 24498
rect 44044 24444 44100 24446
rect 43036 23212 43092 23268
rect 43036 22988 43092 23044
rect 42700 21756 42756 21812
rect 43148 21084 43204 21140
rect 42700 20972 42756 21028
rect 43484 23042 43540 23044
rect 43484 22990 43486 23042
rect 43486 22990 43538 23042
rect 43538 22990 43540 23042
rect 43484 22988 43540 22990
rect 43708 21980 43764 22036
rect 43372 20860 43428 20916
rect 42812 20130 42868 20132
rect 42812 20078 42814 20130
rect 42814 20078 42866 20130
rect 42866 20078 42868 20130
rect 42812 20076 42868 20078
rect 44044 22876 44100 22932
rect 44044 21980 44100 22036
rect 43932 21532 43988 21588
rect 44268 25228 44324 25284
rect 44268 23938 44324 23940
rect 44268 23886 44270 23938
rect 44270 23886 44322 23938
rect 44322 23886 44324 23938
rect 44268 23884 44324 23886
rect 44156 20636 44212 20692
rect 44268 23548 44324 23604
rect 44268 20412 44324 20468
rect 44156 20300 44212 20356
rect 43484 19068 43540 19124
rect 43708 19852 43764 19908
rect 42364 18956 42420 19012
rect 42588 18450 42644 18452
rect 42588 18398 42590 18450
rect 42590 18398 42642 18450
rect 42642 18398 42644 18450
rect 42588 18396 42644 18398
rect 43148 18450 43204 18452
rect 43148 18398 43150 18450
rect 43150 18398 43202 18450
rect 43202 18398 43204 18450
rect 43148 18396 43204 18398
rect 43820 19180 43876 19236
rect 43932 20188 43988 20244
rect 45164 29986 45220 29988
rect 45164 29934 45166 29986
rect 45166 29934 45218 29986
rect 45218 29934 45220 29986
rect 45164 29932 45220 29934
rect 44716 28252 44772 28308
rect 44604 27746 44660 27748
rect 44604 27694 44606 27746
rect 44606 27694 44658 27746
rect 44658 27694 44660 27746
rect 44604 27692 44660 27694
rect 44604 26908 44660 26964
rect 44492 21756 44548 21812
rect 44492 21420 44548 21476
rect 44492 20188 44548 20244
rect 44492 20018 44548 20020
rect 44492 19966 44494 20018
rect 44494 19966 44546 20018
rect 44546 19966 44548 20018
rect 44492 19964 44548 19966
rect 44604 19852 44660 19908
rect 44156 19628 44212 19684
rect 43820 18172 43876 18228
rect 41244 17164 41300 17220
rect 41020 16828 41076 16884
rect 42588 17164 42644 17220
rect 42924 17052 42980 17108
rect 42588 16770 42644 16772
rect 42588 16718 42590 16770
rect 42590 16718 42642 16770
rect 42642 16718 42644 16770
rect 42588 16716 42644 16718
rect 40908 14588 40964 14644
rect 41916 14418 41972 14420
rect 41916 14366 41918 14418
rect 41918 14366 41970 14418
rect 41970 14366 41972 14418
rect 41916 14364 41972 14366
rect 41356 13804 41412 13860
rect 40908 13580 40964 13636
rect 41804 13634 41860 13636
rect 41804 13582 41806 13634
rect 41806 13582 41858 13634
rect 41858 13582 41860 13634
rect 41804 13580 41860 13582
rect 41804 13356 41860 13412
rect 41020 12908 41076 12964
rect 41020 12012 41076 12068
rect 41020 11170 41076 11172
rect 41020 11118 41022 11170
rect 41022 11118 41074 11170
rect 41074 11118 41076 11170
rect 41020 11116 41076 11118
rect 41020 10892 41076 10948
rect 40460 10834 40516 10836
rect 40460 10782 40462 10834
rect 40462 10782 40514 10834
rect 40514 10782 40516 10834
rect 40460 10780 40516 10782
rect 40908 10108 40964 10164
rect 41132 9996 41188 10052
rect 41580 11340 41636 11396
rect 41356 10834 41412 10836
rect 41356 10782 41358 10834
rect 41358 10782 41410 10834
rect 41410 10782 41412 10834
rect 41356 10780 41412 10782
rect 41468 10610 41524 10612
rect 41468 10558 41470 10610
rect 41470 10558 41522 10610
rect 41522 10558 41524 10610
rect 41468 10556 41524 10558
rect 41692 11004 41748 11060
rect 42364 16098 42420 16100
rect 42364 16046 42366 16098
rect 42366 16046 42418 16098
rect 42418 16046 42420 16098
rect 42364 16044 42420 16046
rect 42700 15372 42756 15428
rect 42476 15148 42532 15204
rect 42588 13580 42644 13636
rect 42476 13020 42532 13076
rect 42252 12962 42308 12964
rect 42252 12910 42254 12962
rect 42254 12910 42306 12962
rect 42306 12910 42308 12962
rect 42252 12908 42308 12910
rect 42028 11340 42084 11396
rect 42700 12012 42756 12068
rect 41916 11004 41972 11060
rect 42028 10668 42084 10724
rect 42140 11116 42196 11172
rect 42252 10556 42308 10612
rect 41916 10498 41972 10500
rect 41916 10446 41918 10498
rect 41918 10446 41970 10498
rect 41970 10446 41972 10498
rect 41916 10444 41972 10446
rect 40684 7308 40740 7364
rect 40796 7980 40852 8036
rect 41244 7868 41300 7924
rect 41468 7644 41524 7700
rect 43148 17388 43204 17444
rect 43484 15202 43540 15204
rect 43484 15150 43486 15202
rect 43486 15150 43538 15202
rect 43538 15150 43540 15202
rect 43484 15148 43540 15150
rect 43036 13074 43092 13076
rect 43036 13022 43038 13074
rect 43038 13022 43090 13074
rect 43090 13022 43092 13074
rect 43036 13020 43092 13022
rect 42924 11788 42980 11844
rect 43372 11004 43428 11060
rect 42812 10668 42868 10724
rect 43932 17164 43988 17220
rect 43820 16268 43876 16324
rect 43932 14364 43988 14420
rect 44268 19404 44324 19460
rect 43932 13634 43988 13636
rect 43932 13582 43934 13634
rect 43934 13582 43986 13634
rect 43986 13582 43988 13634
rect 43932 13580 43988 13582
rect 43708 10780 43764 10836
rect 43820 10610 43876 10612
rect 43820 10558 43822 10610
rect 43822 10558 43874 10610
rect 43874 10558 43876 10610
rect 43820 10556 43876 10558
rect 42364 10108 42420 10164
rect 42700 9548 42756 9604
rect 42476 9042 42532 9044
rect 42476 8990 42478 9042
rect 42478 8990 42530 9042
rect 42530 8990 42532 9042
rect 42476 8988 42532 8990
rect 42140 8428 42196 8484
rect 43932 9772 43988 9828
rect 43596 9548 43652 9604
rect 42812 8428 42868 8484
rect 43820 9266 43876 9268
rect 43820 9214 43822 9266
rect 43822 9214 43874 9266
rect 43874 9214 43876 9266
rect 43820 9212 43876 9214
rect 43148 8316 43204 8372
rect 42924 8258 42980 8260
rect 42924 8206 42926 8258
rect 42926 8206 42978 8258
rect 42978 8206 42980 8258
rect 42924 8204 42980 8206
rect 43820 8204 43876 8260
rect 44268 19010 44324 19012
rect 44268 18958 44270 19010
rect 44270 18958 44322 19010
rect 44322 18958 44324 19010
rect 44268 18956 44324 18958
rect 44156 17554 44212 17556
rect 44156 17502 44158 17554
rect 44158 17502 44210 17554
rect 44210 17502 44212 17554
rect 44156 17500 44212 17502
rect 44156 16716 44212 16772
rect 44492 18284 44548 18340
rect 44604 17276 44660 17332
rect 44268 16604 44324 16660
rect 45724 29986 45780 29988
rect 45724 29934 45726 29986
rect 45726 29934 45778 29986
rect 45778 29934 45780 29986
rect 45724 29932 45780 29934
rect 45500 29650 45556 29652
rect 45500 29598 45502 29650
rect 45502 29598 45554 29650
rect 45554 29598 45556 29650
rect 45500 29596 45556 29598
rect 45052 27858 45108 27860
rect 45052 27806 45054 27858
rect 45054 27806 45106 27858
rect 45106 27806 45108 27858
rect 45052 27804 45108 27806
rect 45052 27298 45108 27300
rect 45052 27246 45054 27298
rect 45054 27246 45106 27298
rect 45106 27246 45108 27298
rect 45052 27244 45108 27246
rect 44828 26796 44884 26852
rect 45164 26402 45220 26404
rect 45164 26350 45166 26402
rect 45166 26350 45218 26402
rect 45218 26350 45220 26402
rect 45164 26348 45220 26350
rect 44828 24444 44884 24500
rect 45612 27468 45668 27524
rect 45948 27468 46004 27524
rect 45052 23884 45108 23940
rect 44940 23324 44996 23380
rect 45388 26124 45444 26180
rect 46396 31666 46452 31668
rect 46396 31614 46398 31666
rect 46398 31614 46450 31666
rect 46450 31614 46452 31666
rect 46396 31612 46452 31614
rect 48188 37266 48244 37268
rect 48188 37214 48190 37266
rect 48190 37214 48242 37266
rect 48242 37214 48244 37266
rect 48188 37212 48244 37214
rect 47292 36594 47348 36596
rect 47292 36542 47294 36594
rect 47294 36542 47346 36594
rect 47346 36542 47348 36594
rect 47292 36540 47348 36542
rect 47180 36204 47236 36260
rect 49756 44044 49812 44100
rect 49868 43260 49924 43316
rect 49868 42588 49924 42644
rect 49980 42082 50036 42084
rect 49980 42030 49982 42082
rect 49982 42030 50034 42082
rect 50034 42030 50036 42082
rect 49980 42028 50036 42030
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50876 43708 50932 43764
rect 53228 49868 53284 49924
rect 53228 46562 53284 46564
rect 53228 46510 53230 46562
rect 53230 46510 53282 46562
rect 53282 46510 53284 46562
rect 53228 46508 53284 46510
rect 53004 46172 53060 46228
rect 51100 44716 51156 44772
rect 51996 44940 52052 44996
rect 53228 44994 53284 44996
rect 53228 44942 53230 44994
rect 53230 44942 53282 44994
rect 53282 44942 53284 44994
rect 53228 44940 53284 44942
rect 51324 44098 51380 44100
rect 51324 44046 51326 44098
rect 51326 44046 51378 44098
rect 51378 44046 51380 44098
rect 51324 44044 51380 44046
rect 50652 42642 50708 42644
rect 50652 42590 50654 42642
rect 50654 42590 50706 42642
rect 50706 42590 50708 42642
rect 50652 42588 50708 42590
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50428 42028 50484 42084
rect 50316 41970 50372 41972
rect 50316 41918 50318 41970
rect 50318 41918 50370 41970
rect 50370 41918 50372 41970
rect 50316 41916 50372 41918
rect 49868 39452 49924 39508
rect 49644 39340 49700 39396
rect 49308 37660 49364 37716
rect 49420 37996 49476 38052
rect 48972 37266 49028 37268
rect 48972 37214 48974 37266
rect 48974 37214 49026 37266
rect 49026 37214 49028 37266
rect 48972 37212 49028 37214
rect 48860 35308 48916 35364
rect 48748 34300 48804 34356
rect 49196 35586 49252 35588
rect 49196 35534 49198 35586
rect 49198 35534 49250 35586
rect 49250 35534 49252 35586
rect 49196 35532 49252 35534
rect 49980 39058 50036 39060
rect 49980 39006 49982 39058
rect 49982 39006 50034 39058
rect 50034 39006 50036 39058
rect 49980 39004 50036 39006
rect 49756 37996 49812 38052
rect 49980 38780 50036 38836
rect 49532 37154 49588 37156
rect 49532 37102 49534 37154
rect 49534 37102 49586 37154
rect 49586 37102 49588 37154
rect 49532 37100 49588 37102
rect 49756 36316 49812 36372
rect 49980 35922 50036 35924
rect 49980 35870 49982 35922
rect 49982 35870 50034 35922
rect 50034 35870 50036 35922
rect 49980 35868 50036 35870
rect 50092 36428 50148 36484
rect 49756 35308 49812 35364
rect 48860 34018 48916 34020
rect 48860 33966 48862 34018
rect 48862 33966 48914 34018
rect 48914 33966 48916 34018
rect 48860 33964 48916 33966
rect 47180 33516 47236 33572
rect 47292 33740 47348 33796
rect 47068 29372 47124 29428
rect 48300 29932 48356 29988
rect 48188 29538 48244 29540
rect 48188 29486 48190 29538
rect 48190 29486 48242 29538
rect 48242 29486 48244 29538
rect 48188 29484 48244 29486
rect 47964 29372 48020 29428
rect 47068 28866 47124 28868
rect 47068 28814 47070 28866
rect 47070 28814 47122 28866
rect 47122 28814 47124 28866
rect 47068 28812 47124 28814
rect 46508 28530 46564 28532
rect 46508 28478 46510 28530
rect 46510 28478 46562 28530
rect 46562 28478 46564 28530
rect 46508 28476 46564 28478
rect 47068 27244 47124 27300
rect 46508 27132 46564 27188
rect 47964 28812 48020 28868
rect 48300 28700 48356 28756
rect 46284 24780 46340 24836
rect 46284 23826 46340 23828
rect 46284 23774 46286 23826
rect 46286 23774 46338 23826
rect 46338 23774 46340 23826
rect 46284 23772 46340 23774
rect 45724 23660 45780 23716
rect 45388 23324 45444 23380
rect 45388 22876 45444 22932
rect 45052 21474 45108 21476
rect 45052 21422 45054 21474
rect 45054 21422 45106 21474
rect 45106 21422 45108 21474
rect 45052 21420 45108 21422
rect 45164 20802 45220 20804
rect 45164 20750 45166 20802
rect 45166 20750 45218 20802
rect 45218 20750 45220 20802
rect 45164 20748 45220 20750
rect 45388 20802 45444 20804
rect 45388 20750 45390 20802
rect 45390 20750 45442 20802
rect 45442 20750 45444 20802
rect 45388 20748 45444 20750
rect 44940 20300 44996 20356
rect 45500 20300 45556 20356
rect 45388 20188 45444 20244
rect 45052 20076 45108 20132
rect 44940 19628 44996 19684
rect 44716 16322 44772 16324
rect 44716 16270 44718 16322
rect 44718 16270 44770 16322
rect 44770 16270 44772 16322
rect 44716 16268 44772 16270
rect 44268 16210 44324 16212
rect 44268 16158 44270 16210
rect 44270 16158 44322 16210
rect 44322 16158 44324 16210
rect 44268 16156 44324 16158
rect 44044 8316 44100 8372
rect 42588 8034 42644 8036
rect 42588 7982 42590 8034
rect 42590 7982 42642 8034
rect 42642 7982 42644 8034
rect 42588 7980 42644 7982
rect 42140 7698 42196 7700
rect 42140 7646 42142 7698
rect 42142 7646 42194 7698
rect 42194 7646 42196 7698
rect 42140 7644 42196 7646
rect 41020 7250 41076 7252
rect 41020 7198 41022 7250
rect 41022 7198 41074 7250
rect 41074 7198 41076 7250
rect 41020 7196 41076 7198
rect 41804 7250 41860 7252
rect 41804 7198 41806 7250
rect 41806 7198 41858 7250
rect 41858 7198 41860 7250
rect 41804 7196 41860 7198
rect 43036 7196 43092 7252
rect 42476 6860 42532 6916
rect 44156 14924 44212 14980
rect 43820 6914 43876 6916
rect 43820 6862 43822 6914
rect 43822 6862 43874 6914
rect 43874 6862 43876 6914
rect 43820 6860 43876 6862
rect 40908 5234 40964 5236
rect 40908 5182 40910 5234
rect 40910 5182 40962 5234
rect 40962 5182 40964 5234
rect 40908 5180 40964 5182
rect 41244 4338 41300 4340
rect 41244 4286 41246 4338
rect 41246 4286 41298 4338
rect 41298 4286 41300 4338
rect 41244 4284 41300 4286
rect 43372 6748 43428 6804
rect 43596 6690 43652 6692
rect 43596 6638 43598 6690
rect 43598 6638 43650 6690
rect 43650 6638 43652 6690
rect 43596 6636 43652 6638
rect 44044 6412 44100 6468
rect 42028 4172 42084 4228
rect 43708 4508 43764 4564
rect 41356 3612 41412 3668
rect 42028 3666 42084 3668
rect 42028 3614 42030 3666
rect 42030 3614 42082 3666
rect 42082 3614 42084 3666
rect 42028 3612 42084 3614
rect 44044 4226 44100 4228
rect 44044 4174 44046 4226
rect 44046 4174 44098 4226
rect 44098 4174 44100 4226
rect 44044 4172 44100 4174
rect 43708 3612 43764 3668
rect 35532 3554 35588 3556
rect 35532 3502 35534 3554
rect 35534 3502 35586 3554
rect 35586 3502 35588 3554
rect 35532 3500 35588 3502
rect 35980 3554 36036 3556
rect 35980 3502 35982 3554
rect 35982 3502 36034 3554
rect 36034 3502 36036 3554
rect 35980 3500 36036 3502
rect 38556 3388 38612 3444
rect 39340 3442 39396 3444
rect 39340 3390 39342 3442
rect 39342 3390 39394 3442
rect 39394 3390 39396 3442
rect 39340 3388 39396 3390
rect 39788 3442 39844 3444
rect 39788 3390 39790 3442
rect 39790 3390 39842 3442
rect 39842 3390 39844 3442
rect 39788 3388 39844 3390
rect 43036 3442 43092 3444
rect 43036 3390 43038 3442
rect 43038 3390 43090 3442
rect 43090 3390 43092 3442
rect 43036 3388 43092 3390
rect 45612 20018 45668 20020
rect 45612 19966 45614 20018
rect 45614 19966 45666 20018
rect 45666 19966 45668 20018
rect 45612 19964 45668 19966
rect 45388 19010 45444 19012
rect 45388 18958 45390 19010
rect 45390 18958 45442 19010
rect 45442 18958 45444 19010
rect 45388 18956 45444 18958
rect 45164 17724 45220 17780
rect 44940 17164 44996 17220
rect 45052 16994 45108 16996
rect 45052 16942 45054 16994
rect 45054 16942 45106 16994
rect 45106 16942 45108 16994
rect 45052 16940 45108 16942
rect 44716 14924 44772 14980
rect 45276 15260 45332 15316
rect 45500 17500 45556 17556
rect 45500 16828 45556 16884
rect 45948 20802 46004 20804
rect 45948 20750 45950 20802
rect 45950 20750 46002 20802
rect 46002 20750 46004 20802
rect 45948 20748 46004 20750
rect 46060 19906 46116 19908
rect 46060 19854 46062 19906
rect 46062 19854 46114 19906
rect 46114 19854 46116 19906
rect 46060 19852 46116 19854
rect 45836 19292 45892 19348
rect 45948 17666 46004 17668
rect 45948 17614 45950 17666
rect 45950 17614 46002 17666
rect 46002 17614 46004 17666
rect 45948 17612 46004 17614
rect 45500 15538 45556 15540
rect 45500 15486 45502 15538
rect 45502 15486 45554 15538
rect 45554 15486 45556 15538
rect 45500 15484 45556 15486
rect 45836 15314 45892 15316
rect 45836 15262 45838 15314
rect 45838 15262 45890 15314
rect 45890 15262 45892 15314
rect 45836 15260 45892 15262
rect 45388 14700 45444 14756
rect 45948 14700 46004 14756
rect 45836 14642 45892 14644
rect 45836 14590 45838 14642
rect 45838 14590 45890 14642
rect 45890 14590 45892 14642
rect 45836 14588 45892 14590
rect 44604 13468 44660 13524
rect 44268 6578 44324 6580
rect 44268 6526 44270 6578
rect 44270 6526 44322 6578
rect 44322 6526 44324 6578
rect 44268 6524 44324 6526
rect 44828 11004 44884 11060
rect 44940 11116 44996 11172
rect 45052 10556 45108 10612
rect 45164 11004 45220 11060
rect 45388 13356 45444 13412
rect 45948 13468 46004 13524
rect 45836 13020 45892 13076
rect 46732 23826 46788 23828
rect 46732 23774 46734 23826
rect 46734 23774 46786 23826
rect 46786 23774 46788 23826
rect 46732 23772 46788 23774
rect 46732 21644 46788 21700
rect 46284 20636 46340 20692
rect 46732 20188 46788 20244
rect 46956 25228 47012 25284
rect 48076 28476 48132 28532
rect 48412 27692 48468 27748
rect 47628 27468 47684 27524
rect 47516 27298 47572 27300
rect 47516 27246 47518 27298
rect 47518 27246 47570 27298
rect 47570 27246 47572 27298
rect 47516 27244 47572 27246
rect 47404 23660 47460 23716
rect 47180 22092 47236 22148
rect 48188 24610 48244 24612
rect 48188 24558 48190 24610
rect 48190 24558 48242 24610
rect 48242 24558 48244 24610
rect 48188 24556 48244 24558
rect 47964 22428 48020 22484
rect 47740 21644 47796 21700
rect 46844 20076 46900 20132
rect 47516 20130 47572 20132
rect 47516 20078 47518 20130
rect 47518 20078 47570 20130
rect 47570 20078 47572 20130
rect 47516 20076 47572 20078
rect 47292 20018 47348 20020
rect 47292 19966 47294 20018
rect 47294 19966 47346 20018
rect 47346 19966 47348 20018
rect 47292 19964 47348 19966
rect 46284 18284 46340 18340
rect 47404 17164 47460 17220
rect 46172 15484 46228 15540
rect 46844 16828 46900 16884
rect 46284 15314 46340 15316
rect 46284 15262 46286 15314
rect 46286 15262 46338 15314
rect 46338 15262 46340 15314
rect 46284 15260 46340 15262
rect 46508 15260 46564 15316
rect 46620 16492 46676 16548
rect 46284 14530 46340 14532
rect 46284 14478 46286 14530
rect 46286 14478 46338 14530
rect 46338 14478 46340 14530
rect 46284 14476 46340 14478
rect 45724 12124 45780 12180
rect 45388 10610 45444 10612
rect 45388 10558 45390 10610
rect 45390 10558 45442 10610
rect 45442 10558 45444 10610
rect 45388 10556 45444 10558
rect 45612 11170 45668 11172
rect 45612 11118 45614 11170
rect 45614 11118 45666 11170
rect 45666 11118 45668 11170
rect 45612 11116 45668 11118
rect 46396 13692 46452 13748
rect 45948 11282 46004 11284
rect 45948 11230 45950 11282
rect 45950 11230 46002 11282
rect 46002 11230 46004 11282
rect 45948 11228 46004 11230
rect 46284 11116 46340 11172
rect 47852 19794 47908 19796
rect 47852 19742 47854 19794
rect 47854 19742 47906 19794
rect 47906 19742 47908 19794
rect 47852 19740 47908 19742
rect 48076 20018 48132 20020
rect 48076 19966 48078 20018
rect 48078 19966 48130 20018
rect 48130 19966 48132 20018
rect 48076 19964 48132 19966
rect 47740 19122 47796 19124
rect 47740 19070 47742 19122
rect 47742 19070 47794 19122
rect 47794 19070 47796 19122
rect 47740 19068 47796 19070
rect 47852 17388 47908 17444
rect 47628 15036 47684 15092
rect 47404 14306 47460 14308
rect 47404 14254 47406 14306
rect 47406 14254 47458 14306
rect 47458 14254 47460 14306
rect 47404 14252 47460 14254
rect 46844 13916 46900 13972
rect 46732 13468 46788 13524
rect 48188 13468 48244 13524
rect 46844 11228 46900 11284
rect 46396 10220 46452 10276
rect 46284 10108 46340 10164
rect 44828 6690 44884 6692
rect 44828 6638 44830 6690
rect 44830 6638 44882 6690
rect 44882 6638 44884 6690
rect 44828 6636 44884 6638
rect 44380 5180 44436 5236
rect 44940 5234 44996 5236
rect 44940 5182 44942 5234
rect 44942 5182 44994 5234
rect 44994 5182 44996 5234
rect 44940 5180 44996 5182
rect 45388 9042 45444 9044
rect 45388 8990 45390 9042
rect 45390 8990 45442 9042
rect 45442 8990 45444 9042
rect 45388 8988 45444 8990
rect 45948 9660 46004 9716
rect 46172 9660 46228 9716
rect 45388 7644 45444 7700
rect 46396 9826 46452 9828
rect 46396 9774 46398 9826
rect 46398 9774 46450 9826
rect 46450 9774 46452 9826
rect 46396 9772 46452 9774
rect 47964 10556 48020 10612
rect 47404 10050 47460 10052
rect 47404 9998 47406 10050
rect 47406 9998 47458 10050
rect 47458 9998 47460 10050
rect 47404 9996 47460 9998
rect 47852 9826 47908 9828
rect 47852 9774 47854 9826
rect 47854 9774 47906 9826
rect 47906 9774 47908 9826
rect 47852 9772 47908 9774
rect 45724 6524 45780 6580
rect 47292 8482 47348 8484
rect 47292 8430 47294 8482
rect 47294 8430 47346 8482
rect 47346 8430 47348 8482
rect 47292 8428 47348 8430
rect 46396 6412 46452 6468
rect 46508 8204 46564 8260
rect 47180 8258 47236 8260
rect 47180 8206 47182 8258
rect 47182 8206 47234 8258
rect 47234 8206 47236 8258
rect 47180 8204 47236 8206
rect 46732 7698 46788 7700
rect 46732 7646 46734 7698
rect 46734 7646 46786 7698
rect 46786 7646 46788 7698
rect 46732 7644 46788 7646
rect 47740 7532 47796 7588
rect 46844 7474 46900 7476
rect 46844 7422 46846 7474
rect 46846 7422 46898 7474
rect 46898 7422 46900 7474
rect 46844 7420 46900 7422
rect 48076 9714 48132 9716
rect 48076 9662 48078 9714
rect 48078 9662 48130 9714
rect 48130 9662 48132 9714
rect 48076 9660 48132 9662
rect 48412 23324 48468 23380
rect 48748 33346 48804 33348
rect 48748 33294 48750 33346
rect 48750 33294 48802 33346
rect 48802 33294 48804 33346
rect 48748 33292 48804 33294
rect 49868 35532 49924 35588
rect 49644 34802 49700 34804
rect 49644 34750 49646 34802
rect 49646 34750 49698 34802
rect 49698 34750 49700 34802
rect 49644 34748 49700 34750
rect 49756 34300 49812 34356
rect 49196 33964 49252 34020
rect 49532 33740 49588 33796
rect 49420 33346 49476 33348
rect 49420 33294 49422 33346
rect 49422 33294 49474 33346
rect 49474 33294 49476 33346
rect 49420 33292 49476 33294
rect 49644 33628 49700 33684
rect 50876 41020 50932 41076
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50428 39564 50484 39620
rect 50540 39506 50596 39508
rect 50540 39454 50542 39506
rect 50542 39454 50594 39506
rect 50594 39454 50596 39506
rect 50540 39452 50596 39454
rect 50652 39340 50708 39396
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50428 38834 50484 38836
rect 50428 38782 50430 38834
rect 50430 38782 50482 38834
rect 50482 38782 50484 38834
rect 50428 38780 50484 38782
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50988 36482 51044 36484
rect 50988 36430 50990 36482
rect 50990 36430 51042 36482
rect 51042 36430 51044 36482
rect 50988 36428 51044 36430
rect 53004 43484 53060 43540
rect 53228 42028 53284 42084
rect 51884 40796 51940 40852
rect 53228 39004 53284 39060
rect 53004 38108 53060 38164
rect 51212 36482 51268 36484
rect 51212 36430 51214 36482
rect 51214 36430 51266 36482
rect 51266 36430 51268 36482
rect 51212 36428 51268 36430
rect 50652 36316 50708 36372
rect 50764 36258 50820 36260
rect 50764 36206 50766 36258
rect 50766 36206 50818 36258
rect 50818 36206 50820 36258
rect 50764 36204 50820 36206
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50316 35868 50372 35924
rect 50092 34354 50148 34356
rect 50092 34302 50094 34354
rect 50094 34302 50146 34354
rect 50146 34302 50148 34354
rect 50092 34300 50148 34302
rect 49868 34188 49924 34244
rect 53228 36428 53284 36484
rect 53004 35420 53060 35476
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50204 34018 50260 34020
rect 50204 33966 50206 34018
rect 50206 33966 50258 34018
rect 50258 33966 50260 34018
rect 50204 33964 50260 33966
rect 50092 33852 50148 33908
rect 49084 32450 49140 32452
rect 49084 32398 49086 32450
rect 49086 32398 49138 32450
rect 49138 32398 49140 32450
rect 49084 32396 49140 32398
rect 48860 32338 48916 32340
rect 48860 32286 48862 32338
rect 48862 32286 48914 32338
rect 48914 32286 48916 32338
rect 48860 32284 48916 32286
rect 49868 31554 49924 31556
rect 49868 31502 49870 31554
rect 49870 31502 49922 31554
rect 49922 31502 49924 31554
rect 49868 31500 49924 31502
rect 48972 30828 49028 30884
rect 50652 33740 50708 33796
rect 50876 33964 50932 34020
rect 50988 33122 51044 33124
rect 50988 33070 50990 33122
rect 50990 33070 51042 33122
rect 51042 33070 51044 33122
rect 50988 33068 51044 33070
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 49980 30882 50036 30884
rect 49980 30830 49982 30882
rect 49982 30830 50034 30882
rect 50034 30830 50036 30882
rect 49980 30828 50036 30830
rect 49644 30268 49700 30324
rect 49084 28812 49140 28868
rect 48972 28700 49028 28756
rect 48636 27804 48692 27860
rect 49084 28642 49140 28644
rect 49084 28590 49086 28642
rect 49086 28590 49138 28642
rect 49138 28590 49140 28642
rect 49084 28588 49140 28590
rect 50540 31890 50596 31892
rect 50540 31838 50542 31890
rect 50542 31838 50594 31890
rect 50594 31838 50596 31890
rect 50540 31836 50596 31838
rect 50428 31554 50484 31556
rect 50428 31502 50430 31554
rect 50430 31502 50482 31554
rect 50482 31502 50484 31554
rect 50428 31500 50484 31502
rect 52444 33068 52500 33124
rect 53004 32732 53060 32788
rect 51100 31500 51156 31556
rect 52444 31836 52500 31892
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 49980 29372 50036 29428
rect 49980 27746 50036 27748
rect 49980 27694 49982 27746
rect 49982 27694 50034 27746
rect 50034 27694 50036 27746
rect 49980 27692 50036 27694
rect 52892 30268 52948 30324
rect 48748 24722 48804 24724
rect 48748 24670 48750 24722
rect 48750 24670 48802 24722
rect 48802 24670 48804 24722
rect 48748 24668 48804 24670
rect 48860 24556 48916 24612
rect 48748 23154 48804 23156
rect 48748 23102 48750 23154
rect 48750 23102 48802 23154
rect 48802 23102 48804 23154
rect 48748 23100 48804 23102
rect 48748 19794 48804 19796
rect 48748 19742 48750 19794
rect 48750 19742 48802 19794
rect 48802 19742 48804 19794
rect 48748 19740 48804 19742
rect 48636 18284 48692 18340
rect 48748 18172 48804 18228
rect 49868 26402 49924 26404
rect 49868 26350 49870 26402
rect 49870 26350 49922 26402
rect 49922 26350 49924 26402
rect 49868 26348 49924 26350
rect 49532 25340 49588 25396
rect 49868 26066 49924 26068
rect 49868 26014 49870 26066
rect 49870 26014 49922 26066
rect 49922 26014 49924 26066
rect 49868 26012 49924 26014
rect 49868 25506 49924 25508
rect 49868 25454 49870 25506
rect 49870 25454 49922 25506
rect 49922 25454 49924 25506
rect 49868 25452 49924 25454
rect 49420 24722 49476 24724
rect 49420 24670 49422 24722
rect 49422 24670 49474 24722
rect 49474 24670 49476 24722
rect 49420 24668 49476 24670
rect 49308 23660 49364 23716
rect 49196 23324 49252 23380
rect 49868 24668 49924 24724
rect 49868 23884 49924 23940
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 51212 29538 51268 29540
rect 51212 29486 51214 29538
rect 51214 29486 51266 29538
rect 51266 29486 51268 29538
rect 51212 29484 51268 29486
rect 51884 29426 51940 29428
rect 51884 29374 51886 29426
rect 51886 29374 51938 29426
rect 51938 29374 51940 29426
rect 51884 29372 51940 29374
rect 52444 29426 52500 29428
rect 52444 29374 52446 29426
rect 52446 29374 52498 29426
rect 52498 29374 52500 29426
rect 52444 29372 52500 29374
rect 53228 30098 53284 30100
rect 53228 30046 53230 30098
rect 53230 30046 53282 30098
rect 53282 30046 53284 30098
rect 53228 30044 53284 30046
rect 53116 29372 53172 29428
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 51660 27244 51716 27300
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 52444 27244 52500 27300
rect 53340 27356 53396 27412
rect 52892 26348 52948 26404
rect 50204 25394 50260 25396
rect 50204 25342 50206 25394
rect 50206 25342 50258 25394
rect 50258 25342 50260 25394
rect 50204 25340 50260 25342
rect 50540 25282 50596 25284
rect 50540 25230 50542 25282
rect 50542 25230 50594 25282
rect 50594 25230 50596 25282
rect 50540 25228 50596 25230
rect 51100 25506 51156 25508
rect 51100 25454 51102 25506
rect 51102 25454 51154 25506
rect 51154 25454 51156 25506
rect 51100 25452 51156 25454
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50764 24892 50820 24948
rect 50316 24668 50372 24724
rect 50204 24610 50260 24612
rect 50204 24558 50206 24610
rect 50206 24558 50258 24610
rect 50258 24558 50260 24610
rect 50204 24556 50260 24558
rect 49756 23660 49812 23716
rect 49196 22482 49252 22484
rect 49196 22430 49198 22482
rect 49198 22430 49250 22482
rect 49250 22430 49252 22482
rect 49196 22428 49252 22430
rect 49980 22204 50036 22260
rect 49868 20578 49924 20580
rect 49868 20526 49870 20578
rect 49870 20526 49922 20578
rect 49922 20526 49924 20578
rect 49868 20524 49924 20526
rect 49084 19068 49140 19124
rect 49308 19346 49364 19348
rect 49308 19294 49310 19346
rect 49310 19294 49362 19346
rect 49362 19294 49364 19346
rect 49308 19292 49364 19294
rect 49196 17666 49252 17668
rect 49196 17614 49198 17666
rect 49198 17614 49250 17666
rect 49250 17614 49252 17666
rect 49196 17612 49252 17614
rect 49756 19964 49812 20020
rect 49196 17388 49252 17444
rect 49308 16994 49364 16996
rect 49308 16942 49310 16994
rect 49310 16942 49362 16994
rect 49362 16942 49364 16994
rect 49308 16940 49364 16942
rect 49644 18284 49700 18340
rect 49196 16492 49252 16548
rect 49196 15986 49252 15988
rect 49196 15934 49198 15986
rect 49198 15934 49250 15986
rect 49250 15934 49252 15986
rect 49196 15932 49252 15934
rect 49084 15484 49140 15540
rect 49084 15314 49140 15316
rect 49084 15262 49086 15314
rect 49086 15262 49138 15314
rect 49138 15262 49140 15314
rect 49084 15260 49140 15262
rect 48636 15148 48692 15204
rect 48524 14252 48580 14308
rect 49196 13468 49252 13524
rect 49756 15986 49812 15988
rect 49756 15934 49758 15986
rect 49758 15934 49810 15986
rect 49810 15934 49812 15986
rect 49756 15932 49812 15934
rect 49980 15986 50036 15988
rect 49980 15934 49982 15986
rect 49982 15934 50034 15986
rect 50034 15934 50036 15986
rect 49980 15932 50036 15934
rect 49644 15484 49700 15540
rect 50092 15372 50148 15428
rect 49084 12124 49140 12180
rect 48300 9212 48356 9268
rect 48188 8204 48244 8260
rect 48300 7532 48356 7588
rect 45164 4956 45220 5012
rect 44492 4562 44548 4564
rect 44492 4510 44494 4562
rect 44494 4510 44546 4562
rect 44546 4510 44548 4562
rect 44492 4508 44548 4510
rect 46732 6636 46788 6692
rect 47404 6690 47460 6692
rect 47404 6638 47406 6690
rect 47406 6638 47458 6690
rect 47458 6638 47460 6690
rect 47404 6636 47460 6638
rect 47628 6690 47684 6692
rect 47628 6638 47630 6690
rect 47630 6638 47682 6690
rect 47682 6638 47684 6690
rect 47628 6636 47684 6638
rect 47180 6578 47236 6580
rect 47180 6526 47182 6578
rect 47182 6526 47234 6578
rect 47234 6526 47236 6578
rect 47180 6524 47236 6526
rect 46732 5122 46788 5124
rect 46732 5070 46734 5122
rect 46734 5070 46786 5122
rect 46786 5070 46788 5122
rect 46732 5068 46788 5070
rect 48076 6690 48132 6692
rect 48076 6638 48078 6690
rect 48078 6638 48130 6690
rect 48130 6638 48132 6690
rect 48076 6636 48132 6638
rect 49196 11116 49252 11172
rect 49196 10108 49252 10164
rect 49084 9660 49140 9716
rect 48412 6972 48468 7028
rect 48524 7420 48580 7476
rect 50876 24834 50932 24836
rect 50876 24782 50878 24834
rect 50878 24782 50930 24834
rect 50930 24782 50932 24834
rect 50876 24780 50932 24782
rect 50428 23938 50484 23940
rect 50428 23886 50430 23938
rect 50430 23886 50482 23938
rect 50482 23886 50484 23938
rect 50428 23884 50484 23886
rect 51324 25116 51380 25172
rect 51660 26012 51716 26068
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50876 23100 50932 23156
rect 50988 22258 51044 22260
rect 50988 22206 50990 22258
rect 50990 22206 51042 22258
rect 51042 22206 51044 22258
rect 50988 22204 51044 22206
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50316 20188 50372 20244
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50316 19292 50372 19348
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 51436 22258 51492 22260
rect 51436 22206 51438 22258
rect 51438 22206 51490 22258
rect 51490 22206 51492 22258
rect 51436 22204 51492 22206
rect 51660 24722 51716 24724
rect 51660 24670 51662 24722
rect 51662 24670 51714 24722
rect 51714 24670 51716 24722
rect 51660 24668 51716 24670
rect 52108 23772 52164 23828
rect 51324 19852 51380 19908
rect 53228 24722 53284 24724
rect 53228 24670 53230 24722
rect 53230 24670 53282 24722
rect 53282 24670 53284 24722
rect 53228 24668 53284 24670
rect 52892 23660 52948 23716
rect 53116 23154 53172 23156
rect 53116 23102 53118 23154
rect 53118 23102 53170 23154
rect 53170 23102 53172 23154
rect 53116 23100 53172 23102
rect 52668 22258 52724 22260
rect 52668 22206 52670 22258
rect 52670 22206 52722 22258
rect 52722 22206 52724 22258
rect 52668 22204 52724 22206
rect 53228 21980 53284 22036
rect 52668 21698 52724 21700
rect 52668 21646 52670 21698
rect 52670 21646 52722 21698
rect 52722 21646 52724 21698
rect 52668 21644 52724 21646
rect 51548 20524 51604 20580
rect 51772 19852 51828 19908
rect 50988 18396 51044 18452
rect 51212 17948 51268 18004
rect 52220 19346 52276 19348
rect 52220 19294 52222 19346
rect 52222 19294 52274 19346
rect 52274 19294 52276 19346
rect 52220 19292 52276 19294
rect 51884 18450 51940 18452
rect 51884 18398 51886 18450
rect 51886 18398 51938 18450
rect 51938 18398 51940 18450
rect 51884 18396 51940 18398
rect 52444 18450 52500 18452
rect 52444 18398 52446 18450
rect 52446 18398 52498 18450
rect 52498 18398 52500 18450
rect 52444 18396 52500 18398
rect 52220 18172 52276 18228
rect 51772 17948 51828 18004
rect 52108 17948 52164 18004
rect 50988 17612 51044 17668
rect 51212 17612 51268 17668
rect 50652 17554 50708 17556
rect 50652 17502 50654 17554
rect 50654 17502 50706 17554
rect 50706 17502 50708 17554
rect 50652 17500 50708 17502
rect 50540 17388 50596 17444
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 51100 17388 51156 17444
rect 50876 16380 50932 16436
rect 51324 17106 51380 17108
rect 51324 17054 51326 17106
rect 51326 17054 51378 17106
rect 51378 17054 51380 17106
rect 51324 17052 51380 17054
rect 51884 17388 51940 17444
rect 51772 17106 51828 17108
rect 51772 17054 51774 17106
rect 51774 17054 51826 17106
rect 51826 17054 51828 17106
rect 51772 17052 51828 17054
rect 51548 16604 51604 16660
rect 50428 15986 50484 15988
rect 50428 15934 50430 15986
rect 50430 15934 50482 15986
rect 50482 15934 50484 15986
rect 50428 15932 50484 15934
rect 50652 15874 50708 15876
rect 50652 15822 50654 15874
rect 50654 15822 50706 15874
rect 50706 15822 50708 15874
rect 50652 15820 50708 15822
rect 51324 15820 51380 15876
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50316 15484 50372 15540
rect 51100 15314 51156 15316
rect 51100 15262 51102 15314
rect 51102 15262 51154 15314
rect 51154 15262 51156 15314
rect 51100 15260 51156 15262
rect 51324 15202 51380 15204
rect 51324 15150 51326 15202
rect 51326 15150 51378 15202
rect 51378 15150 51380 15202
rect 51324 15148 51380 15150
rect 50204 14588 50260 14644
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 51100 13468 51156 13524
rect 50316 13356 50372 13412
rect 49532 12178 49588 12180
rect 49532 12126 49534 12178
rect 49534 12126 49586 12178
rect 49586 12126 49588 12178
rect 49532 12124 49588 12126
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 51436 13356 51492 13412
rect 49532 11170 49588 11172
rect 49532 11118 49534 11170
rect 49534 11118 49586 11170
rect 49586 11118 49588 11170
rect 49532 11116 49588 11118
rect 49420 10610 49476 10612
rect 49420 10558 49422 10610
rect 49422 10558 49474 10610
rect 49474 10558 49476 10610
rect 49420 10556 49476 10558
rect 49644 10834 49700 10836
rect 49644 10782 49646 10834
rect 49646 10782 49698 10834
rect 49698 10782 49700 10834
rect 49644 10780 49700 10782
rect 50652 11116 50708 11172
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 49756 9772 49812 9828
rect 49868 9714 49924 9716
rect 49868 9662 49870 9714
rect 49870 9662 49922 9714
rect 49922 9662 49924 9714
rect 49868 9660 49924 9662
rect 49756 8988 49812 9044
rect 49196 6972 49252 7028
rect 48636 6636 48692 6692
rect 47852 6412 47908 6468
rect 49532 6578 49588 6580
rect 49532 6526 49534 6578
rect 49534 6526 49586 6578
rect 49586 6526 49588 6578
rect 49532 6524 49588 6526
rect 48860 5068 48916 5124
rect 50092 9548 50148 9604
rect 50204 7532 50260 7588
rect 49980 6748 50036 6804
rect 50204 6412 50260 6468
rect 50540 9714 50596 9716
rect 50540 9662 50542 9714
rect 50542 9662 50594 9714
rect 50594 9662 50596 9714
rect 50540 9660 50596 9662
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50428 7532 50484 7588
rect 51772 15820 51828 15876
rect 52780 17500 52836 17556
rect 52556 17388 52612 17444
rect 53228 21698 53284 21700
rect 53228 21646 53230 21698
rect 53230 21646 53282 21698
rect 53282 21646 53284 21698
rect 53228 21644 53284 21646
rect 53228 19906 53284 19908
rect 53228 19854 53230 19906
rect 53230 19854 53282 19906
rect 53282 19854 53284 19906
rect 53228 19852 53284 19854
rect 53228 19292 53284 19348
rect 53004 17612 53060 17668
rect 52892 16994 52948 16996
rect 52892 16942 52894 16994
rect 52894 16942 52946 16994
rect 52946 16942 52948 16994
rect 52892 16940 52948 16942
rect 52668 16882 52724 16884
rect 52668 16830 52670 16882
rect 52670 16830 52722 16882
rect 52722 16830 52724 16882
rect 52668 16828 52724 16830
rect 53228 16882 53284 16884
rect 53228 16830 53230 16882
rect 53230 16830 53282 16882
rect 53282 16830 53284 16882
rect 53228 16828 53284 16830
rect 52668 15986 52724 15988
rect 52668 15934 52670 15986
rect 52670 15934 52722 15986
rect 52722 15934 52724 15986
rect 52668 15932 52724 15934
rect 52780 15874 52836 15876
rect 52780 15822 52782 15874
rect 52782 15822 52834 15874
rect 52834 15822 52836 15874
rect 52780 15820 52836 15822
rect 52332 15538 52388 15540
rect 52332 15486 52334 15538
rect 52334 15486 52386 15538
rect 52386 15486 52388 15538
rect 52332 15484 52388 15486
rect 53116 15372 53172 15428
rect 52108 15202 52164 15204
rect 52108 15150 52110 15202
rect 52110 15150 52162 15202
rect 52162 15150 52164 15202
rect 52108 15148 52164 15150
rect 52668 15036 52724 15092
rect 52220 13468 52276 13524
rect 52668 14364 52724 14420
rect 51996 12012 52052 12068
rect 52220 11282 52276 11284
rect 52220 11230 52222 11282
rect 52222 11230 52274 11282
rect 52274 11230 52276 11282
rect 52220 11228 52276 11230
rect 52220 9042 52276 9044
rect 52220 8990 52222 9042
rect 52222 8990 52274 9042
rect 52274 8990 52276 9042
rect 52220 8988 52276 8990
rect 52332 7586 52388 7588
rect 52332 7534 52334 7586
rect 52334 7534 52386 7586
rect 52386 7534 52388 7586
rect 52332 7532 52388 7534
rect 52892 14252 52948 14308
rect 53340 13970 53396 13972
rect 53340 13918 53342 13970
rect 53342 13918 53394 13970
rect 53394 13918 53396 13970
rect 53340 13916 53396 13918
rect 53228 12066 53284 12068
rect 53228 12014 53230 12066
rect 53230 12014 53282 12066
rect 53282 12014 53284 12066
rect 53228 12012 53284 12014
rect 53228 11282 53284 11284
rect 53228 11230 53230 11282
rect 53230 11230 53282 11282
rect 53282 11230 53284 11282
rect 53228 11228 53284 11230
rect 52780 9660 52836 9716
rect 53228 8540 53284 8596
rect 51548 6636 51604 6692
rect 52668 6690 52724 6692
rect 52668 6638 52670 6690
rect 52670 6638 52722 6690
rect 52722 6638 52724 6690
rect 52668 6636 52724 6638
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 52220 6466 52276 6468
rect 52220 6414 52222 6466
rect 52222 6414 52274 6466
rect 52274 6414 52276 6466
rect 52220 6412 52276 6414
rect 53228 6466 53284 6468
rect 53228 6414 53230 6466
rect 53230 6414 53282 6466
rect 53282 6414 53284 6466
rect 53228 6412 53284 6414
rect 53340 5852 53396 5908
rect 49980 5122 50036 5124
rect 49980 5070 49982 5122
rect 49982 5070 50034 5122
rect 50034 5070 50036 5122
rect 49980 5068 50036 5070
rect 49980 4450 50036 4452
rect 49980 4398 49982 4450
rect 49982 4398 50034 4450
rect 50034 4398 50036 4450
rect 49980 4396 50036 4398
rect 52668 4956 52724 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 51100 4450 51156 4452
rect 51100 4398 51102 4450
rect 51102 4398 51154 4450
rect 51154 4398 51156 4450
rect 51100 4396 51156 4398
rect 50652 3836 50708 3892
rect 49644 3666 49700 3668
rect 49644 3614 49646 3666
rect 49646 3614 49698 3666
rect 49698 3614 49700 3666
rect 49644 3612 49700 3614
rect 44156 3388 44212 3444
rect 47404 3442 47460 3444
rect 47404 3390 47406 3442
rect 47406 3390 47458 3442
rect 47458 3390 47460 3442
rect 47404 3388 47460 3390
rect 51996 3612 52052 3668
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 53228 3836 53284 3892
rect 52444 3164 52500 3220
rect 53228 3164 53284 3220
<< metal3 >>
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 54200 51604 55000 51632
rect 51090 51548 51100 51604
rect 51156 51548 55000 51604
rect 54200 51520 55000 51548
rect 49858 51324 49868 51380
rect 49924 51324 51660 51380
rect 51716 51324 51726 51380
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 23090 50652 23100 50708
rect 23156 50652 26124 50708
rect 26180 50652 26190 50708
rect 26338 50652 26348 50708
rect 26404 50652 31276 50708
rect 31332 50652 31342 50708
rect 16930 50540 16940 50596
rect 16996 50540 17948 50596
rect 18004 50540 20188 50596
rect 20244 50540 20254 50596
rect 32386 50540 32396 50596
rect 32452 50540 35756 50596
rect 35812 50540 35822 50596
rect 39890 50540 39900 50596
rect 39956 50540 42700 50596
rect 42756 50540 43036 50596
rect 43092 50540 43372 50596
rect 43428 50540 45724 50596
rect 45780 50540 45790 50596
rect 49186 50540 49196 50596
rect 49252 50540 49756 50596
rect 49812 50540 51436 50596
rect 51492 50540 51502 50596
rect 17602 50428 17612 50484
rect 17668 50428 21420 50484
rect 21476 50428 21486 50484
rect 21830 50428 21868 50484
rect 21924 50428 21934 50484
rect 22082 50428 22092 50484
rect 22148 50428 22988 50484
rect 23044 50428 23436 50484
rect 23492 50428 23996 50484
rect 24052 50428 24062 50484
rect 24322 50428 24332 50484
rect 24388 50428 26012 50484
rect 26068 50428 29148 50484
rect 29204 50428 29214 50484
rect 33170 50428 33180 50484
rect 33236 50428 33964 50484
rect 34020 50428 34030 50484
rect 37650 50428 37660 50484
rect 37716 50428 39116 50484
rect 39172 50428 39182 50484
rect 41010 50428 41020 50484
rect 41076 50428 42364 50484
rect 42420 50428 42430 50484
rect 49970 50428 49980 50484
rect 50036 50428 51212 50484
rect 51268 50428 51278 50484
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 19618 49980 19628 50036
rect 19684 49980 20412 50036
rect 20468 49980 21196 50036
rect 21252 49980 21262 50036
rect 35074 49980 35084 50036
rect 35140 49980 36764 50036
rect 36820 49980 36830 50036
rect 37202 49980 37212 50036
rect 37268 49980 39788 50036
rect 39844 49980 39854 50036
rect 19842 49868 19852 49924
rect 19908 49868 23324 49924
rect 23380 49868 23390 49924
rect 25890 49868 25900 49924
rect 25956 49868 27356 49924
rect 27412 49868 27422 49924
rect 33842 49868 33852 49924
rect 33908 49868 37772 49924
rect 37828 49868 41132 49924
rect 41188 49868 42028 49924
rect 42084 49868 42094 49924
rect 42354 49868 42364 49924
rect 42420 49868 43484 49924
rect 43540 49868 43550 49924
rect 48962 49868 48972 49924
rect 49028 49868 53228 49924
rect 53284 49868 53294 49924
rect 21298 49756 21308 49812
rect 21364 49756 22988 49812
rect 23044 49756 23548 49812
rect 23604 49756 23614 49812
rect 26786 49756 26796 49812
rect 26852 49756 27692 49812
rect 27748 49756 27758 49812
rect 34402 49756 34412 49812
rect 34468 49756 34748 49812
rect 34804 49756 36652 49812
rect 36708 49756 39004 49812
rect 39060 49756 39070 49812
rect 46050 49756 46060 49812
rect 46116 49756 48860 49812
rect 48916 49756 48926 49812
rect 26562 49644 26572 49700
rect 26628 49644 31388 49700
rect 31444 49644 31454 49700
rect 36866 49644 36876 49700
rect 36932 49644 37548 49700
rect 37604 49644 37614 49700
rect 39890 49644 39900 49700
rect 39956 49644 40908 49700
rect 40964 49644 40974 49700
rect 20066 49532 20076 49588
rect 20132 49532 21644 49588
rect 21700 49532 21710 49588
rect 28018 49532 28028 49588
rect 28084 49532 29260 49588
rect 29316 49532 29326 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 22428 49196 26348 49252
rect 26404 49196 26414 49252
rect 20738 48972 20748 49028
rect 20804 48972 21756 49028
rect 21812 48972 21822 49028
rect 22428 48916 22484 49196
rect 23622 49084 23660 49140
rect 23716 49084 25564 49140
rect 25620 49084 25630 49140
rect 23538 48972 23548 49028
rect 23604 48972 25788 49028
rect 25844 48972 25854 49028
rect 54200 48916 55000 48944
rect 22418 48860 22428 48916
rect 22484 48860 22494 48916
rect 23986 48860 23996 48916
rect 24052 48860 24556 48916
rect 24612 48860 25340 48916
rect 25396 48860 27132 48916
rect 27188 48860 37772 48916
rect 37828 48860 37838 48916
rect 39778 48860 39788 48916
rect 39844 48860 41132 48916
rect 41188 48860 41198 48916
rect 42242 48860 42252 48916
rect 42308 48860 42700 48916
rect 42756 48860 42766 48916
rect 51874 48860 51884 48916
rect 51940 48860 55000 48916
rect 54200 48832 55000 48860
rect 22306 48748 22316 48804
rect 22372 48748 22876 48804
rect 22932 48748 24108 48804
rect 24164 48748 24444 48804
rect 24500 48748 24510 48804
rect 26674 48748 26684 48804
rect 26740 48748 27468 48804
rect 27524 48748 27534 48804
rect 33954 48748 33964 48804
rect 34020 48748 35084 48804
rect 35140 48748 35150 48804
rect 42018 48748 42028 48804
rect 42084 48748 42476 48804
rect 42532 48748 42542 48804
rect 46610 48748 46620 48804
rect 46676 48748 47180 48804
rect 47236 48748 47246 48804
rect 23538 48636 23548 48692
rect 23604 48636 23642 48692
rect 34850 48636 34860 48692
rect 34916 48636 36988 48692
rect 37044 48636 37054 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 47170 48300 47180 48356
rect 47236 48300 48972 48356
rect 49028 48300 49038 48356
rect 23622 48188 23660 48244
rect 23716 48188 23726 48244
rect 34290 48188 34300 48244
rect 34356 48188 34972 48244
rect 35028 48188 35038 48244
rect 33394 48076 33404 48132
rect 33460 48076 34524 48132
rect 34580 48076 34590 48132
rect 46498 48076 46508 48132
rect 46564 48076 47404 48132
rect 47460 48076 48188 48132
rect 48244 48076 49196 48132
rect 49252 48076 49262 48132
rect 46610 47964 46620 48020
rect 46676 47964 47740 48020
rect 47796 47964 47806 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 22754 47628 22764 47684
rect 22820 47628 27916 47684
rect 27972 47628 27982 47684
rect 37762 47628 37772 47684
rect 37828 47628 39228 47684
rect 39284 47628 42364 47684
rect 42420 47628 43148 47684
rect 43204 47628 43214 47684
rect 49074 47516 49084 47572
rect 49140 47516 49644 47572
rect 49700 47516 49710 47572
rect 13010 47404 13020 47460
rect 13076 47404 16268 47460
rect 16324 47404 17948 47460
rect 18004 47404 18014 47460
rect 20514 47404 20524 47460
rect 20580 47404 22428 47460
rect 22484 47404 22494 47460
rect 40226 47404 40236 47460
rect 40292 47404 42588 47460
rect 42644 47404 45500 47460
rect 45556 47404 45566 47460
rect 47730 47404 47740 47460
rect 47796 47404 49532 47460
rect 49588 47404 49598 47460
rect 16930 47292 16940 47348
rect 16996 47292 21420 47348
rect 21476 47292 21486 47348
rect 21830 47292 21868 47348
rect 21924 47292 25900 47348
rect 25956 47292 26908 47348
rect 26964 47292 26974 47348
rect 31938 47292 31948 47348
rect 32004 47292 35196 47348
rect 35252 47292 35262 47348
rect 26114 47180 26124 47236
rect 26180 47180 28252 47236
rect 28308 47180 31164 47236
rect 31220 47180 33180 47236
rect 33236 47180 33246 47236
rect 37314 47180 37324 47236
rect 37380 47180 39228 47236
rect 39284 47180 39294 47236
rect 42028 47180 42812 47236
rect 42868 47180 42878 47236
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 42028 47012 42084 47180
rect 40002 46956 40012 47012
rect 40068 46956 41804 47012
rect 41860 46956 42084 47012
rect 43652 47068 45948 47124
rect 46004 47068 46014 47124
rect 43652 46900 43708 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 17938 46844 17948 46900
rect 18004 46844 19292 46900
rect 19348 46844 19358 46900
rect 26898 46844 26908 46900
rect 26964 46844 43708 46900
rect 19618 46732 19628 46788
rect 19684 46732 20524 46788
rect 20580 46732 21084 46788
rect 21140 46732 21150 46788
rect 28018 46732 28028 46788
rect 28084 46732 30044 46788
rect 30100 46732 30110 46788
rect 40348 46732 41580 46788
rect 41636 46732 41646 46788
rect 41794 46732 41804 46788
rect 41860 46732 42588 46788
rect 42644 46732 42654 46788
rect 40348 46676 40404 46732
rect 15810 46620 15820 46676
rect 15876 46620 16380 46676
rect 16436 46620 17500 46676
rect 17556 46620 18732 46676
rect 18788 46620 18798 46676
rect 20626 46620 20636 46676
rect 20692 46620 22764 46676
rect 22820 46620 23212 46676
rect 23268 46620 23278 46676
rect 36866 46620 36876 46676
rect 36932 46620 39900 46676
rect 39956 46620 40348 46676
rect 40404 46620 40414 46676
rect 41234 46620 41244 46676
rect 41300 46620 42924 46676
rect 42980 46620 42990 46676
rect 43362 46620 43372 46676
rect 43428 46620 45276 46676
rect 45332 46620 50428 46676
rect 50484 46620 50494 46676
rect 13682 46508 13692 46564
rect 13748 46508 16268 46564
rect 16324 46508 16334 46564
rect 41804 46452 41860 46620
rect 43026 46508 43036 46564
rect 43092 46508 44156 46564
rect 44212 46508 44222 46564
rect 48850 46508 48860 46564
rect 48916 46508 53228 46564
rect 53284 46508 53294 46564
rect 41794 46396 41804 46452
rect 41860 46396 41870 46452
rect 38882 46284 38892 46340
rect 38948 46284 45836 46340
rect 45892 46284 47740 46340
rect 47796 46284 48748 46340
rect 48804 46284 48814 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 54200 46228 55000 46256
rect 36418 46172 36428 46228
rect 36484 46172 37660 46228
rect 37716 46172 37726 46228
rect 52994 46172 53004 46228
rect 53060 46172 55000 46228
rect 54200 46144 55000 46172
rect 20290 46060 20300 46116
rect 20356 46060 21644 46116
rect 21700 46060 23100 46116
rect 23156 46060 23166 46116
rect 48290 45948 48300 46004
rect 48356 45948 49196 46004
rect 49252 45948 49262 46004
rect 16930 45836 16940 45892
rect 16996 45836 17948 45892
rect 18004 45836 22988 45892
rect 23044 45836 23054 45892
rect 24770 45836 24780 45892
rect 24836 45836 25900 45892
rect 25956 45836 27804 45892
rect 27860 45836 27870 45892
rect 42802 45836 42812 45892
rect 42868 45836 43708 45892
rect 10434 45724 10444 45780
rect 10500 45724 11228 45780
rect 11284 45724 11294 45780
rect 13906 45724 13916 45780
rect 13972 45724 14812 45780
rect 14868 45724 17612 45780
rect 17668 45724 18508 45780
rect 18564 45724 24108 45780
rect 24164 45724 24668 45780
rect 24724 45724 24734 45780
rect 35970 45724 35980 45780
rect 36036 45724 37324 45780
rect 37380 45724 37884 45780
rect 37940 45724 37950 45780
rect 43652 45668 43708 45836
rect 15922 45612 15932 45668
rect 15988 45612 16268 45668
rect 16324 45612 16334 45668
rect 23538 45612 23548 45668
rect 23604 45612 24444 45668
rect 24500 45612 24510 45668
rect 25330 45612 25340 45668
rect 25396 45612 26348 45668
rect 26404 45612 26414 45668
rect 43652 45612 46284 45668
rect 46340 45612 46350 45668
rect 43652 45500 49084 45556
rect 49140 45500 49150 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 7298 45388 7308 45444
rect 7364 45388 9772 45444
rect 9828 45388 9838 45444
rect 43652 45332 43708 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 11106 45276 11116 45332
rect 11172 45276 12348 45332
rect 12404 45276 12414 45332
rect 21970 45276 21980 45332
rect 22036 45276 22988 45332
rect 23044 45276 23054 45332
rect 24658 45276 24668 45332
rect 24724 45276 33124 45332
rect 40002 45276 40012 45332
rect 40068 45276 43708 45332
rect 43810 45276 43820 45332
rect 43876 45276 44268 45332
rect 44324 45276 46620 45332
rect 46676 45276 46686 45332
rect 47842 45276 47852 45332
rect 47908 45276 48748 45332
rect 48804 45276 48814 45332
rect 33068 45220 33124 45276
rect 12226 45164 12236 45220
rect 12292 45164 12684 45220
rect 12740 45164 12908 45220
rect 12964 45164 12974 45220
rect 20066 45164 20076 45220
rect 20132 45164 22316 45220
rect 22372 45164 22652 45220
rect 22708 45164 28812 45220
rect 28868 45164 28878 45220
rect 33058 45164 33068 45220
rect 33124 45164 33134 45220
rect 42354 45164 42364 45220
rect 42420 45164 44156 45220
rect 44212 45164 44222 45220
rect 12450 45052 12460 45108
rect 12516 45052 14252 45108
rect 14308 45052 14318 45108
rect 17826 45052 17836 45108
rect 17892 45052 19516 45108
rect 19572 45052 19582 45108
rect 25666 45052 25676 45108
rect 25732 45052 29260 45108
rect 29316 45052 29596 45108
rect 29652 45052 30716 45108
rect 30772 45052 30782 45108
rect 32386 45052 32396 45108
rect 32452 45052 33852 45108
rect 33908 45052 35308 45108
rect 35364 45052 36092 45108
rect 36148 45052 36158 45108
rect 37090 45052 37100 45108
rect 37156 45052 38220 45108
rect 38276 45052 38780 45108
rect 38836 45052 38846 45108
rect 41906 45052 41916 45108
rect 41972 45052 42476 45108
rect 42532 45052 42542 45108
rect 11554 44940 11564 44996
rect 11620 44940 12572 44996
rect 12628 44940 12638 44996
rect 22418 44940 22428 44996
rect 22484 44940 25116 44996
rect 25172 44940 25182 44996
rect 25778 44940 25788 44996
rect 25844 44940 28140 44996
rect 28196 44940 28206 44996
rect 34850 44940 34860 44996
rect 34916 44940 37212 44996
rect 37268 44940 43708 44996
rect 43764 44940 43774 44996
rect 51100 44940 51996 44996
rect 52052 44940 53228 44996
rect 53284 44940 53294 44996
rect 12572 44884 12628 44940
rect 12572 44828 12796 44884
rect 12852 44828 12862 44884
rect 19842 44828 19852 44884
rect 19908 44828 23996 44884
rect 24052 44828 24062 44884
rect 33506 44828 33516 44884
rect 33572 44828 47068 44884
rect 47124 44828 47516 44884
rect 47572 44828 47582 44884
rect 51100 44772 51156 44940
rect 19730 44716 19740 44772
rect 19796 44716 21980 44772
rect 22036 44716 22316 44772
rect 22372 44716 22382 44772
rect 51090 44716 51100 44772
rect 51156 44716 51166 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 10882 44492 10892 44548
rect 10948 44492 11788 44548
rect 11844 44492 12908 44548
rect 12964 44492 12974 44548
rect 22866 44492 22876 44548
rect 22932 44492 25900 44548
rect 25956 44492 25966 44548
rect 32050 44492 32060 44548
rect 32116 44492 33852 44548
rect 33908 44492 34188 44548
rect 34244 44492 34748 44548
rect 34804 44492 35532 44548
rect 35588 44492 35598 44548
rect 9650 44380 9660 44436
rect 9716 44380 10444 44436
rect 10500 44380 10510 44436
rect 11890 44380 11900 44436
rect 11956 44380 12572 44436
rect 12628 44380 13356 44436
rect 13412 44380 22092 44436
rect 22148 44380 22158 44436
rect 31938 44380 31948 44436
rect 32004 44380 32732 44436
rect 32788 44380 32798 44436
rect 35074 44380 35084 44436
rect 35140 44380 37100 44436
rect 37156 44380 37166 44436
rect 11330 44268 11340 44324
rect 11396 44268 12684 44324
rect 12740 44268 12750 44324
rect 17266 44268 17276 44324
rect 17332 44268 17724 44324
rect 17780 44268 19292 44324
rect 19348 44268 19358 44324
rect 32386 44268 32396 44324
rect 32452 44268 33628 44324
rect 33684 44268 33694 44324
rect 38546 44268 38556 44324
rect 38612 44268 39004 44324
rect 39060 44268 39452 44324
rect 39508 44268 39518 44324
rect 40674 44268 40684 44324
rect 40740 44268 41132 44324
rect 41188 44268 45052 44324
rect 45108 44268 45612 44324
rect 45668 44268 45678 44324
rect 12786 44156 12796 44212
rect 12852 44156 13580 44212
rect 13636 44156 14140 44212
rect 14196 44156 14206 44212
rect 14466 44156 14476 44212
rect 14532 44156 15148 44212
rect 15204 44156 15932 44212
rect 15988 44156 16828 44212
rect 16884 44156 16894 44212
rect 33506 44156 33516 44212
rect 33572 44156 34636 44212
rect 34692 44156 35756 44212
rect 35812 44156 37772 44212
rect 37828 44156 37838 44212
rect 44258 44156 44268 44212
rect 44324 44156 44940 44212
rect 44996 44156 45006 44212
rect 9650 44044 9660 44100
rect 9716 44044 10780 44100
rect 10836 44044 10846 44100
rect 16482 44044 16492 44100
rect 16548 44044 17388 44100
rect 17444 44044 17454 44100
rect 39778 44044 39788 44100
rect 39844 44044 40348 44100
rect 40404 44044 40414 44100
rect 49746 44044 49756 44100
rect 49812 44044 51324 44100
rect 51380 44044 51390 44100
rect 10882 43932 10892 43988
rect 10948 43932 14700 43988
rect 14756 43932 17948 43988
rect 18004 43932 18014 43988
rect 36082 43932 36092 43988
rect 36148 43932 38780 43988
rect 38836 43932 38846 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 9986 43820 9996 43876
rect 10052 43820 11452 43876
rect 11508 43820 11518 43876
rect 12002 43820 12012 43876
rect 12068 43820 17500 43876
rect 17556 43820 17566 43876
rect 34178 43820 34188 43876
rect 34244 43820 37884 43876
rect 37940 43820 37950 43876
rect 17500 43764 17556 43820
rect 17500 43708 19068 43764
rect 19124 43708 20076 43764
rect 20132 43708 20142 43764
rect 36306 43708 36316 43764
rect 36372 43708 39452 43764
rect 39508 43708 40012 43764
rect 40068 43708 40078 43764
rect 43698 43708 43708 43764
rect 43764 43708 50876 43764
rect 50932 43708 50942 43764
rect 7522 43596 7532 43652
rect 7588 43596 9772 43652
rect 9828 43596 9838 43652
rect 16146 43596 16156 43652
rect 16212 43596 19404 43652
rect 19460 43596 19470 43652
rect 22642 43596 22652 43652
rect 22708 43596 24108 43652
rect 24164 43596 24174 43652
rect 26114 43596 26124 43652
rect 26180 43596 26572 43652
rect 26628 43596 26638 43652
rect 28354 43596 28364 43652
rect 28420 43596 28812 43652
rect 28868 43596 34412 43652
rect 34468 43596 34478 43652
rect 41346 43596 41356 43652
rect 41412 43596 43484 43652
rect 43540 43596 44492 43652
rect 44548 43596 45388 43652
rect 45444 43596 46060 43652
rect 46116 43596 46732 43652
rect 46788 43596 46798 43652
rect 54200 43540 55000 43568
rect 10882 43484 10892 43540
rect 10948 43484 11788 43540
rect 11844 43484 11854 43540
rect 41458 43484 41468 43540
rect 41524 43484 42588 43540
rect 42644 43484 42654 43540
rect 52994 43484 53004 43540
rect 53060 43484 55000 43540
rect 32162 43372 32172 43428
rect 32228 43372 35980 43428
rect 36036 43372 36046 43428
rect 38612 43372 39788 43428
rect 39844 43372 39854 43428
rect 38612 43316 38668 43372
rect 15474 43260 15484 43316
rect 15540 43260 16828 43316
rect 16884 43260 16894 43316
rect 18946 43260 18956 43316
rect 19012 43260 31500 43316
rect 31556 43260 32060 43316
rect 32116 43260 32126 43316
rect 32386 43260 32396 43316
rect 32452 43260 38668 43316
rect 19730 43148 19740 43204
rect 19796 43148 20412 43204
rect 20468 43148 22764 43204
rect 22820 43148 34188 43204
rect 34244 43148 34254 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 42588 43092 42644 43484
rect 54200 43456 55000 43484
rect 48850 43260 48860 43316
rect 48916 43260 49868 43316
rect 49924 43260 49934 43316
rect 16706 43036 16716 43092
rect 16772 43036 17612 43092
rect 17668 43036 21980 43092
rect 22036 43036 22046 43092
rect 42588 43036 48524 43092
rect 48580 43036 48590 43092
rect 17042 42924 17052 42980
rect 17108 42924 28364 42980
rect 28420 42924 28430 42980
rect 31378 42924 31388 42980
rect 31444 42924 31724 42980
rect 31780 42924 41132 42980
rect 41188 42924 41468 42980
rect 41524 42924 41534 42980
rect 25442 42812 25452 42868
rect 25508 42812 26348 42868
rect 26404 42812 26414 42868
rect 26674 42812 26684 42868
rect 26740 42812 27020 42868
rect 27076 42812 27086 42868
rect 32050 42812 32060 42868
rect 32116 42812 32732 42868
rect 32788 42812 32798 42868
rect 19170 42700 19180 42756
rect 19236 42700 21308 42756
rect 21364 42700 21374 42756
rect 23650 42700 23660 42756
rect 23716 42700 25004 42756
rect 25060 42700 25340 42756
rect 25396 42700 25406 42756
rect 26852 42700 27916 42756
rect 27972 42700 29260 42756
rect 29316 42700 29326 42756
rect 29698 42700 29708 42756
rect 29764 42700 34524 42756
rect 34580 42700 34590 42756
rect 38546 42700 38556 42756
rect 38612 42700 40348 42756
rect 40404 42700 40414 42756
rect 47058 42700 47068 42756
rect 47124 42700 47404 42756
rect 47460 42700 47470 42756
rect 23874 42588 23884 42644
rect 23940 42588 24444 42644
rect 24500 42588 25228 42644
rect 25284 42588 25294 42644
rect 14802 42476 14812 42532
rect 14868 42476 18060 42532
rect 18116 42476 18126 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 26852 42308 26908 42700
rect 35074 42588 35084 42644
rect 35140 42588 35980 42644
rect 36036 42588 36046 42644
rect 49858 42588 49868 42644
rect 49924 42588 50652 42644
rect 50708 42588 50718 42644
rect 27458 42476 27468 42532
rect 27524 42476 28588 42532
rect 28644 42476 29484 42532
rect 29540 42476 29550 42532
rect 33618 42476 33628 42532
rect 33684 42476 34412 42532
rect 34468 42476 34478 42532
rect 35858 42476 35868 42532
rect 35924 42476 38220 42532
rect 38276 42476 38286 42532
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 15092 42252 19684 42308
rect 21970 42252 21980 42308
rect 22036 42252 22428 42308
rect 22484 42252 26908 42308
rect 36978 42252 36988 42308
rect 37044 42252 41916 42308
rect 41972 42252 41982 42308
rect 15092 42196 15148 42252
rect 19628 42196 19684 42252
rect 11666 42140 11676 42196
rect 11732 42140 15148 42196
rect 16034 42140 16044 42196
rect 16100 42140 16110 42196
rect 19628 42140 25788 42196
rect 25844 42140 25854 42196
rect 12226 42028 12236 42084
rect 12292 42028 13020 42084
rect 13076 42028 13086 42084
rect 16044 41972 16100 42140
rect 25788 42084 25844 42140
rect 25788 42028 26124 42084
rect 26180 42028 27468 42084
rect 27524 42028 27534 42084
rect 34514 42028 34524 42084
rect 34580 42028 35084 42084
rect 35140 42028 35868 42084
rect 35924 42028 35934 42084
rect 44930 42028 44940 42084
rect 44996 42028 46284 42084
rect 46340 42028 46350 42084
rect 49970 42028 49980 42084
rect 50036 42028 50428 42084
rect 50484 42028 53228 42084
rect 53284 42028 53294 42084
rect 10434 41916 10444 41972
rect 10500 41916 12908 41972
rect 12964 41916 12974 41972
rect 13682 41916 13692 41972
rect 13748 41916 16100 41972
rect 21522 41916 21532 41972
rect 21588 41916 23212 41972
rect 23268 41916 24556 41972
rect 24612 41916 25116 41972
rect 25172 41916 25182 41972
rect 26338 41916 26348 41972
rect 26404 41916 29820 41972
rect 29876 41916 30380 41972
rect 30436 41916 30446 41972
rect 37090 41916 37100 41972
rect 37156 41916 41020 41972
rect 41076 41916 41086 41972
rect 47954 41916 47964 41972
rect 48020 41916 49084 41972
rect 49140 41916 50316 41972
rect 50372 41916 50382 41972
rect 8082 41804 8092 41860
rect 8148 41804 10556 41860
rect 10612 41804 10622 41860
rect 21746 41804 21756 41860
rect 21812 41804 24220 41860
rect 24276 41804 29148 41860
rect 29204 41804 29214 41860
rect 29362 41804 29372 41860
rect 29428 41804 31948 41860
rect 32004 41804 32014 41860
rect 45042 41804 45052 41860
rect 45108 41804 46732 41860
rect 46788 41804 46798 41860
rect 20402 41692 20412 41748
rect 20468 41692 21308 41748
rect 21364 41692 23100 41748
rect 23156 41692 23996 41748
rect 24052 41692 24062 41748
rect 34066 41692 34076 41748
rect 34132 41692 34972 41748
rect 35028 41692 35038 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 17938 41244 17948 41300
rect 18004 41244 20636 41300
rect 20692 41244 20702 41300
rect 33618 41244 33628 41300
rect 33684 41244 38108 41300
rect 38164 41244 38556 41300
rect 38612 41244 38622 41300
rect 40114 41244 40124 41300
rect 40180 41244 42588 41300
rect 42644 41244 43484 41300
rect 43540 41244 43550 41300
rect 10210 41132 10220 41188
rect 10276 41132 10892 41188
rect 10948 41132 10958 41188
rect 12674 41132 12684 41188
rect 12740 41132 13692 41188
rect 13748 41132 13758 41188
rect 18722 41132 18732 41188
rect 18788 41132 19628 41188
rect 19684 41132 19694 41188
rect 20514 41132 20524 41188
rect 20580 41132 22652 41188
rect 22708 41132 22718 41188
rect 36194 41132 36204 41188
rect 36260 41132 37212 41188
rect 37268 41132 37278 41188
rect 11106 41020 11116 41076
rect 11172 41020 12124 41076
rect 12180 41020 12572 41076
rect 12628 41020 12908 41076
rect 12964 41020 12974 41076
rect 18050 41020 18060 41076
rect 18116 41020 18508 41076
rect 18564 41020 18574 41076
rect 18946 41020 18956 41076
rect 19012 41020 20188 41076
rect 20244 41020 21196 41076
rect 21252 41020 21262 41076
rect 31042 41020 31052 41076
rect 31108 41020 33852 41076
rect 33908 41020 33918 41076
rect 34290 41020 34300 41076
rect 34356 41020 37100 41076
rect 37156 41020 37166 41076
rect 49186 41020 49196 41076
rect 49252 41020 50876 41076
rect 50932 41020 50942 41076
rect 16146 40908 16156 40964
rect 16212 40908 18620 40964
rect 18676 40908 18686 40964
rect 36642 40908 36652 40964
rect 36708 40908 37324 40964
rect 37380 40908 37390 40964
rect 43138 40908 43148 40964
rect 43204 40908 44156 40964
rect 44212 40908 44222 40964
rect 54200 40852 55000 40880
rect 51874 40796 51884 40852
rect 51940 40796 55000 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 54200 40768 55000 40796
rect 20514 40684 20524 40740
rect 20580 40684 21532 40740
rect 21588 40684 21598 40740
rect 38546 40684 38556 40740
rect 38612 40684 39452 40740
rect 39508 40684 43708 40740
rect 10770 40572 10780 40628
rect 10836 40572 11228 40628
rect 11284 40572 30044 40628
rect 30100 40572 30110 40628
rect 30706 40572 30716 40628
rect 30772 40572 34300 40628
rect 34356 40572 34366 40628
rect 39666 40572 39676 40628
rect 39732 40572 40124 40628
rect 40180 40572 40908 40628
rect 40964 40572 40974 40628
rect 43652 40516 43708 40684
rect 30594 40460 30604 40516
rect 30660 40460 33964 40516
rect 34020 40460 34030 40516
rect 41906 40460 41916 40516
rect 41972 40460 43036 40516
rect 43092 40460 43102 40516
rect 43652 40460 43932 40516
rect 43988 40460 43998 40516
rect 10882 40348 10892 40404
rect 10948 40348 11900 40404
rect 11956 40348 11966 40404
rect 17826 40348 17836 40404
rect 17892 40348 18396 40404
rect 18452 40348 19068 40404
rect 19124 40348 22428 40404
rect 22484 40348 22494 40404
rect 29810 40348 29820 40404
rect 29876 40348 33180 40404
rect 33236 40348 33246 40404
rect 42018 40348 42028 40404
rect 42084 40348 44044 40404
rect 44100 40348 44110 40404
rect 42028 40292 42084 40348
rect 37986 40236 37996 40292
rect 38052 40236 38780 40292
rect 38836 40236 38846 40292
rect 41234 40236 41244 40292
rect 41300 40236 42084 40292
rect 45154 40236 45164 40292
rect 45220 40236 48524 40292
rect 48580 40236 48590 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 13794 39788 13804 39844
rect 13860 39788 14140 39844
rect 14196 39788 14206 39844
rect 26852 39788 36988 39844
rect 37044 39788 37054 39844
rect 8372 39676 8988 39732
rect 9044 39676 11564 39732
rect 11620 39676 11630 39732
rect 15474 39676 15484 39732
rect 15540 39676 17500 39732
rect 17556 39676 17836 39732
rect 17892 39676 18172 39732
rect 18228 39676 18956 39732
rect 19012 39676 21644 39732
rect 21700 39676 22092 39732
rect 22148 39676 22158 39732
rect 8372 39620 8428 39676
rect 5730 39564 5740 39620
rect 5796 39564 7308 39620
rect 7364 39564 8428 39620
rect 10098 39452 10108 39508
rect 10164 39452 11228 39508
rect 11284 39452 11294 39508
rect 15484 39396 15540 39676
rect 26852 39620 26908 39788
rect 12114 39340 12124 39396
rect 12180 39340 15540 39396
rect 15596 39564 26908 39620
rect 27682 39564 27692 39620
rect 27748 39564 28364 39620
rect 28420 39564 29260 39620
rect 29316 39564 29326 39620
rect 33506 39564 33516 39620
rect 33572 39564 34188 39620
rect 34244 39564 34254 39620
rect 49186 39564 49196 39620
rect 49252 39564 50428 39620
rect 50484 39564 50494 39620
rect 15596 39284 15652 39564
rect 44034 39452 44044 39508
rect 44100 39452 44828 39508
rect 44884 39452 44894 39508
rect 49858 39452 49868 39508
rect 49924 39452 50540 39508
rect 50596 39452 50606 39508
rect 18946 39340 18956 39396
rect 19012 39340 25340 39396
rect 25396 39340 25406 39396
rect 32498 39340 32508 39396
rect 32564 39340 33628 39396
rect 33684 39340 33694 39396
rect 49634 39340 49644 39396
rect 49700 39340 50652 39396
rect 50708 39340 50718 39396
rect 12002 39228 12012 39284
rect 12068 39228 15652 39284
rect 20962 39228 20972 39284
rect 21028 39228 22092 39284
rect 22148 39228 22158 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 38770 39116 38780 39172
rect 38836 39116 39340 39172
rect 39396 39116 39406 39172
rect 44930 39116 44940 39172
rect 44996 39116 46396 39172
rect 46452 39116 46462 39172
rect 10994 39004 11004 39060
rect 11060 39004 11676 39060
rect 11732 39004 25452 39060
rect 25508 39004 30716 39060
rect 30772 39004 30782 39060
rect 43698 39004 43708 39060
rect 43764 39004 44380 39060
rect 44436 39004 44446 39060
rect 8372 38892 9772 38948
rect 9828 38892 9838 38948
rect 12786 38892 12796 38948
rect 12852 38892 13916 38948
rect 13972 38892 13982 38948
rect 8372 38836 8428 38892
rect 44940 38836 44996 39116
rect 49970 39004 49980 39060
rect 50036 39004 53228 39060
rect 53284 39004 53294 39060
rect 6514 38780 6524 38836
rect 6580 38780 8428 38836
rect 38098 38780 38108 38836
rect 38164 38780 41356 38836
rect 41412 38780 43708 38836
rect 43810 38780 43820 38836
rect 43876 38780 44996 38836
rect 49970 38780 49980 38836
rect 50036 38780 50428 38836
rect 50484 38780 50494 38836
rect 43652 38724 43708 38780
rect 29362 38668 29372 38724
rect 29428 38668 37212 38724
rect 37268 38668 38220 38724
rect 38276 38668 38286 38724
rect 43652 38668 44044 38724
rect 44100 38668 45500 38724
rect 45556 38668 45566 38724
rect 27010 38556 27020 38612
rect 27076 38556 28476 38612
rect 28532 38556 36036 38612
rect 35980 38500 36036 38556
rect 35970 38444 35980 38500
rect 36036 38444 36046 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 27906 38332 27916 38388
rect 27972 38332 29820 38388
rect 29876 38332 29886 38388
rect 28578 38220 28588 38276
rect 28644 38220 29708 38276
rect 29764 38220 29774 38276
rect 54200 38164 55000 38192
rect 33506 38108 33516 38164
rect 33572 38108 35532 38164
rect 35588 38108 37100 38164
rect 37156 38108 38556 38164
rect 38612 38108 38622 38164
rect 52994 38108 53004 38164
rect 53060 38108 55000 38164
rect 54200 38080 55000 38108
rect 28578 37996 28588 38052
rect 28644 37996 29484 38052
rect 29540 37996 29550 38052
rect 49410 37996 49420 38052
rect 49476 37996 49756 38052
rect 49812 37996 49822 38052
rect 16370 37884 16380 37940
rect 16436 37884 46060 37940
rect 46116 37884 46126 37940
rect 6850 37772 6860 37828
rect 6916 37772 7532 37828
rect 7588 37772 7598 37828
rect 16706 37772 16716 37828
rect 16772 37772 27020 37828
rect 27076 37772 27086 37828
rect 44370 37660 44380 37716
rect 44436 37660 49308 37716
rect 49364 37660 49374 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 25666 37436 25676 37492
rect 25732 37436 29036 37492
rect 29092 37436 29102 37492
rect 18162 37324 18172 37380
rect 18228 37324 19628 37380
rect 19684 37324 19694 37380
rect 26114 37324 26124 37380
rect 26180 37324 30828 37380
rect 30884 37324 30894 37380
rect 5282 37212 5292 37268
rect 5348 37212 6748 37268
rect 6804 37212 6814 37268
rect 17938 37212 17948 37268
rect 18004 37212 18844 37268
rect 18900 37212 18910 37268
rect 48178 37212 48188 37268
rect 48244 37212 48972 37268
rect 49028 37212 49038 37268
rect 2482 37100 2492 37156
rect 2548 37100 5740 37156
rect 5796 37100 5806 37156
rect 6850 37100 6860 37156
rect 6916 37100 6926 37156
rect 7522 37100 7532 37156
rect 7588 37100 8540 37156
rect 8596 37100 9884 37156
rect 9940 37100 9950 37156
rect 18274 37100 18284 37156
rect 18340 37100 19852 37156
rect 19908 37100 19918 37156
rect 45154 37100 45164 37156
rect 45220 37100 45836 37156
rect 45892 37100 45902 37156
rect 46162 37100 46172 37156
rect 46228 37100 49532 37156
rect 49588 37100 49598 37156
rect 6860 36932 6916 37100
rect 6860 36876 9548 36932
rect 9604 36876 9614 36932
rect 11778 36876 11788 36932
rect 11844 36876 17836 36932
rect 17892 36876 17902 36932
rect 39218 36876 39228 36932
rect 39284 36876 40236 36932
rect 40292 36876 40302 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 14130 36764 14140 36820
rect 14196 36764 18172 36820
rect 18228 36764 18238 36820
rect 15474 36652 15484 36708
rect 15540 36652 16492 36708
rect 16548 36652 16558 36708
rect 45714 36540 45724 36596
rect 45780 36540 47292 36596
rect 47348 36540 47358 36596
rect 22866 36428 22876 36484
rect 22932 36428 25340 36484
rect 25396 36428 25406 36484
rect 39106 36428 39116 36484
rect 39172 36428 40572 36484
rect 40628 36428 43036 36484
rect 43092 36428 43708 36484
rect 43764 36428 44828 36484
rect 44884 36428 44894 36484
rect 50082 36428 50092 36484
rect 50148 36428 50988 36484
rect 51044 36428 51054 36484
rect 51202 36428 51212 36484
rect 51268 36428 53228 36484
rect 53284 36428 53294 36484
rect 22642 36316 22652 36372
rect 22708 36316 24332 36372
rect 24388 36316 24398 36372
rect 31826 36316 31836 36372
rect 31892 36316 45948 36372
rect 46004 36316 46014 36372
rect 49746 36316 49756 36372
rect 49812 36316 50652 36372
rect 50708 36316 50718 36372
rect 6290 36204 6300 36260
rect 6356 36204 9212 36260
rect 9268 36204 9278 36260
rect 9986 36204 9996 36260
rect 10052 36204 10668 36260
rect 10724 36204 10734 36260
rect 30146 36204 30156 36260
rect 30212 36204 38332 36260
rect 38388 36204 38892 36260
rect 38948 36204 38958 36260
rect 44258 36204 44268 36260
rect 44324 36204 45164 36260
rect 45220 36204 45230 36260
rect 47170 36204 47180 36260
rect 47236 36204 50764 36260
rect 50820 36204 50830 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 5730 35868 5740 35924
rect 5796 35868 6636 35924
rect 6692 35868 6702 35924
rect 9986 35868 9996 35924
rect 10052 35868 11788 35924
rect 11844 35868 11854 35924
rect 16034 35868 16044 35924
rect 16100 35868 16604 35924
rect 16660 35868 27132 35924
rect 27188 35868 27198 35924
rect 32610 35868 32620 35924
rect 32676 35868 40236 35924
rect 40292 35868 40302 35924
rect 49970 35868 49980 35924
rect 50036 35868 50316 35924
rect 50372 35868 50382 35924
rect 9538 35756 9548 35812
rect 9604 35756 12460 35812
rect 12516 35756 12526 35812
rect 41234 35756 41244 35812
rect 41300 35756 42924 35812
rect 42980 35756 44268 35812
rect 44324 35756 44828 35812
rect 44884 35756 44894 35812
rect 5058 35644 5068 35700
rect 5124 35644 6524 35700
rect 6580 35644 9772 35700
rect 9828 35644 15596 35700
rect 15652 35644 15662 35700
rect 19730 35644 19740 35700
rect 19796 35644 20412 35700
rect 20468 35644 20478 35700
rect 25778 35644 25788 35700
rect 25844 35644 26348 35700
rect 26404 35644 26796 35700
rect 26852 35644 26862 35700
rect 31602 35644 31612 35700
rect 31668 35644 32284 35700
rect 32340 35644 33180 35700
rect 33236 35644 33246 35700
rect 35522 35644 35532 35700
rect 35588 35644 38892 35700
rect 38948 35644 38958 35700
rect 39442 35644 39452 35700
rect 39508 35644 42140 35700
rect 42196 35644 42206 35700
rect 13346 35532 13356 35588
rect 13412 35532 14028 35588
rect 14084 35532 16716 35588
rect 16772 35532 16782 35588
rect 29474 35532 29484 35588
rect 29540 35532 30156 35588
rect 30212 35532 30222 35588
rect 34626 35532 34636 35588
rect 34692 35532 38220 35588
rect 38276 35532 38286 35588
rect 44146 35532 44156 35588
rect 44212 35532 45276 35588
rect 45332 35532 45342 35588
rect 49186 35532 49196 35588
rect 49252 35532 49868 35588
rect 49924 35532 49934 35588
rect 54200 35476 55000 35504
rect 10658 35420 10668 35476
rect 10724 35420 12012 35476
rect 12068 35420 12796 35476
rect 12852 35420 12862 35476
rect 16930 35420 16940 35476
rect 16996 35420 23100 35476
rect 23156 35420 24220 35476
rect 24276 35420 24286 35476
rect 35186 35420 35196 35476
rect 35252 35420 36092 35476
rect 36148 35420 36158 35476
rect 42802 35420 42812 35476
rect 42868 35420 43596 35476
rect 43652 35420 43662 35476
rect 52994 35420 53004 35476
rect 53060 35420 55000 35476
rect 54200 35392 55000 35420
rect 12114 35308 12124 35364
rect 12180 35308 12460 35364
rect 12516 35308 25340 35364
rect 25396 35308 27132 35364
rect 27188 35308 34076 35364
rect 34132 35308 34636 35364
rect 34692 35308 34702 35364
rect 40114 35308 40124 35364
rect 40180 35308 43708 35364
rect 43764 35308 43774 35364
rect 43922 35308 43932 35364
rect 43988 35308 43998 35364
rect 48850 35308 48860 35364
rect 48916 35308 49756 35364
rect 49812 35308 49822 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 43932 35252 43988 35308
rect 21970 35196 21980 35252
rect 22036 35196 23436 35252
rect 23492 35196 23502 35252
rect 38612 35196 38780 35252
rect 38836 35196 38846 35252
rect 43362 35196 43372 35252
rect 43428 35196 43988 35252
rect 33506 35084 33516 35140
rect 33572 35084 35980 35140
rect 36036 35084 37884 35140
rect 37940 35084 37950 35140
rect 38612 35028 38668 35196
rect 38994 35084 39004 35140
rect 39060 35084 43708 35140
rect 43764 35084 43774 35140
rect 1810 34972 1820 35028
rect 1876 34972 4844 35028
rect 4900 34972 5180 35028
rect 5236 34972 8428 35028
rect 8484 34972 8988 35028
rect 9044 34972 9054 35028
rect 17490 34972 17500 35028
rect 17556 34972 20524 35028
rect 20580 34972 20590 35028
rect 24210 34972 24220 35028
rect 24276 34972 29484 35028
rect 29540 34972 30156 35028
rect 30212 34972 31052 35028
rect 31108 34972 31118 35028
rect 31276 34972 37436 35028
rect 37492 34972 38668 35028
rect 38770 34972 38780 35028
rect 38836 34972 39228 35028
rect 39284 34972 39294 35028
rect 45154 34972 45164 35028
rect 45220 34972 46732 35028
rect 46788 34972 46798 35028
rect 31276 34916 31332 34972
rect 9202 34860 9212 34916
rect 9268 34860 10332 34916
rect 10388 34860 10398 34916
rect 30594 34860 30604 34916
rect 30660 34860 31276 34916
rect 31332 34860 31342 34916
rect 32386 34860 32396 34916
rect 32452 34860 33404 34916
rect 33460 34860 38668 34916
rect 39106 34860 39116 34916
rect 39172 34860 39788 34916
rect 39844 34860 39854 34916
rect 40002 34860 40012 34916
rect 40068 34860 40106 34916
rect 40226 34860 40236 34916
rect 40292 34860 45276 34916
rect 45332 34860 45342 34916
rect 38612 34804 38668 34860
rect 2482 34748 2492 34804
rect 2548 34748 6524 34804
rect 6580 34748 6590 34804
rect 24658 34748 24668 34804
rect 24724 34748 25676 34804
rect 25732 34748 25742 34804
rect 29026 34748 29036 34804
rect 29092 34748 29708 34804
rect 29764 34748 30940 34804
rect 30996 34748 31948 34804
rect 32004 34748 32014 34804
rect 34290 34748 34300 34804
rect 34356 34748 35532 34804
rect 35588 34748 35598 34804
rect 38612 34748 41580 34804
rect 41636 34748 42252 34804
rect 42308 34748 42476 34804
rect 42532 34748 42542 34804
rect 45602 34748 45612 34804
rect 45668 34748 49644 34804
rect 49700 34748 49710 34804
rect 7522 34636 7532 34692
rect 7588 34636 9660 34692
rect 9716 34636 11004 34692
rect 11060 34636 15708 34692
rect 15764 34636 18172 34692
rect 18228 34636 18238 34692
rect 29922 34636 29932 34692
rect 29988 34636 30604 34692
rect 30660 34636 32620 34692
rect 32676 34636 32686 34692
rect 38546 34636 38556 34692
rect 38612 34636 38780 34692
rect 38836 34636 38846 34692
rect 38994 34636 39004 34692
rect 39060 34636 39070 34692
rect 40226 34636 40236 34692
rect 40292 34636 40302 34692
rect 44370 34636 44380 34692
rect 44436 34636 45052 34692
rect 45108 34636 45118 34692
rect 39004 34580 39060 34636
rect 38434 34524 38444 34580
rect 38500 34524 39060 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 6178 34412 6188 34468
rect 6244 34412 8092 34468
rect 8148 34412 8158 34468
rect 11890 34412 11900 34468
rect 11956 34412 18620 34468
rect 18676 34412 18686 34468
rect 34514 34412 34524 34468
rect 34580 34412 35420 34468
rect 35476 34412 37212 34468
rect 37268 34412 39564 34468
rect 39620 34412 40012 34468
rect 40068 34412 40078 34468
rect 40236 34356 40292 34636
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 7522 34300 7532 34356
rect 7588 34300 7868 34356
rect 7924 34300 10444 34356
rect 10500 34300 10510 34356
rect 34178 34300 34188 34356
rect 34244 34300 34860 34356
rect 34916 34300 35196 34356
rect 35252 34300 35980 34356
rect 36036 34300 36046 34356
rect 37874 34300 37884 34356
rect 37940 34300 38668 34356
rect 38770 34300 38780 34356
rect 38836 34300 40292 34356
rect 44370 34300 44380 34356
rect 44436 34300 48748 34356
rect 48804 34300 48814 34356
rect 49746 34300 49756 34356
rect 49812 34300 50092 34356
rect 50148 34300 50158 34356
rect 6738 34188 6748 34244
rect 6804 34188 7196 34244
rect 7252 34188 7262 34244
rect 12226 34188 12236 34244
rect 12292 34188 13580 34244
rect 13636 34188 13646 34244
rect 22418 34188 22428 34244
rect 22484 34188 24332 34244
rect 24388 34188 24398 34244
rect 33282 34188 33292 34244
rect 33348 34188 33964 34244
rect 34020 34188 34030 34244
rect 34962 34188 34972 34244
rect 35028 34188 35756 34244
rect 35812 34188 35822 34244
rect 38612 34188 38668 34300
rect 38724 34188 38734 34244
rect 49858 34188 49868 34244
rect 49924 34188 49934 34244
rect 4610 34076 4620 34132
rect 4676 34076 5292 34132
rect 5348 34076 7420 34132
rect 7476 34076 8988 34132
rect 9044 34076 12012 34132
rect 12068 34076 12078 34132
rect 12674 34076 12684 34132
rect 12740 34076 15036 34132
rect 15092 34076 15102 34132
rect 34514 34076 34524 34132
rect 34580 34076 35868 34132
rect 35924 34076 35934 34132
rect 38546 34076 38556 34132
rect 38612 34076 44156 34132
rect 44212 34076 44222 34132
rect 12562 33964 12572 34020
rect 12628 33964 12908 34020
rect 12964 33964 21980 34020
rect 22036 33964 26908 34020
rect 27122 33964 27132 34020
rect 27188 33964 28252 34020
rect 28308 33964 30604 34020
rect 30660 33964 32396 34020
rect 32452 33964 32462 34020
rect 41570 33964 41580 34020
rect 41636 33964 42588 34020
rect 42644 33964 42924 34020
rect 42980 33964 42990 34020
rect 48850 33964 48860 34020
rect 48916 33964 49196 34020
rect 49252 33964 49262 34020
rect 9650 33852 9660 33908
rect 9716 33852 10052 33908
rect 8978 33740 8988 33796
rect 9044 33740 9548 33796
rect 9604 33740 9614 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 6962 33628 6972 33684
rect 7028 33628 9660 33684
rect 9716 33628 9726 33684
rect 9996 33572 10052 33852
rect 26852 33684 26908 33964
rect 49868 33908 49924 34188
rect 50194 33964 50204 34020
rect 50260 33964 50876 34020
rect 50932 33964 50942 34020
rect 33506 33852 33516 33908
rect 33572 33852 34412 33908
rect 34468 33852 34478 33908
rect 49868 33852 50092 33908
rect 50148 33852 50158 33908
rect 45042 33740 45052 33796
rect 45108 33740 47292 33796
rect 47348 33740 47358 33796
rect 49522 33740 49532 33796
rect 49588 33740 50652 33796
rect 50708 33740 50718 33796
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 26852 33628 31892 33684
rect 37538 33628 37548 33684
rect 37604 33628 38444 33684
rect 38500 33628 38510 33684
rect 42578 33628 42588 33684
rect 42644 33628 49644 33684
rect 49700 33628 49710 33684
rect 31836 33572 31892 33628
rect 8866 33516 8876 33572
rect 8932 33516 9772 33572
rect 9828 33516 9838 33572
rect 9996 33516 11228 33572
rect 11284 33516 11294 33572
rect 31836 33516 33740 33572
rect 33796 33516 33806 33572
rect 43474 33516 43484 33572
rect 43540 33516 47180 33572
rect 47236 33516 47246 33572
rect 9996 33460 10052 33516
rect 5730 33404 5740 33460
rect 5796 33404 7980 33460
rect 8036 33404 10052 33460
rect 16258 33404 16268 33460
rect 16324 33404 24892 33460
rect 24948 33404 25564 33460
rect 25620 33404 25630 33460
rect 32386 33404 32396 33460
rect 32452 33404 32844 33460
rect 32900 33404 33964 33460
rect 34020 33404 35644 33460
rect 35700 33404 37436 33460
rect 37492 33404 37502 33460
rect 24770 33292 24780 33348
rect 24836 33292 41692 33348
rect 41748 33292 42028 33348
rect 42084 33292 42094 33348
rect 44482 33292 44492 33348
rect 44548 33292 45388 33348
rect 45444 33292 46060 33348
rect 46116 33292 48748 33348
rect 48804 33292 49420 33348
rect 49476 33292 49486 33348
rect 26226 33180 26236 33236
rect 26292 33180 27020 33236
rect 27076 33180 27086 33236
rect 37090 33180 37100 33236
rect 37156 33180 38668 33236
rect 38612 33124 38668 33180
rect 10210 33068 10220 33124
rect 10276 33068 11004 33124
rect 11060 33068 11788 33124
rect 11844 33068 11854 33124
rect 14466 33068 14476 33124
rect 14532 33068 15484 33124
rect 15540 33068 15550 33124
rect 17378 33068 17388 33124
rect 17444 33068 17948 33124
rect 18004 33068 31164 33124
rect 31220 33068 31230 33124
rect 37202 33068 37212 33124
rect 37268 33068 38108 33124
rect 38164 33068 38174 33124
rect 38612 33068 41244 33124
rect 41300 33068 41310 33124
rect 42130 33068 42140 33124
rect 42196 33068 42476 33124
rect 42532 33068 43036 33124
rect 43092 33068 45052 33124
rect 45108 33068 45724 33124
rect 45780 33068 45790 33124
rect 50978 33068 50988 33124
rect 51044 33068 52444 33124
rect 52500 33068 52510 33124
rect 26852 32956 41580 33012
rect 41636 32956 41646 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 26852 32900 26908 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 24322 32844 24332 32900
rect 24388 32844 26908 32900
rect 39218 32844 39228 32900
rect 39284 32844 43148 32900
rect 43204 32844 43214 32900
rect 54200 32788 55000 32816
rect 33506 32732 33516 32788
rect 33572 32732 36988 32788
rect 37044 32732 38668 32788
rect 38724 32732 39116 32788
rect 39172 32732 39182 32788
rect 52994 32732 53004 32788
rect 53060 32732 55000 32788
rect 54200 32704 55000 32732
rect 14914 32620 14924 32676
rect 14980 32620 15484 32676
rect 15540 32620 15550 32676
rect 37762 32620 37772 32676
rect 37828 32620 38668 32676
rect 38612 32564 38668 32620
rect 4946 32508 4956 32564
rect 5012 32508 5628 32564
rect 5684 32508 5694 32564
rect 21970 32508 21980 32564
rect 22036 32508 22652 32564
rect 22708 32508 25452 32564
rect 25508 32508 26348 32564
rect 26404 32508 26414 32564
rect 38612 32508 41804 32564
rect 41860 32508 41870 32564
rect 43250 32508 43260 32564
rect 43316 32508 44156 32564
rect 44212 32508 44222 32564
rect 44930 32508 44940 32564
rect 44996 32508 45612 32564
rect 45668 32508 45678 32564
rect 1810 32396 1820 32452
rect 1876 32396 5180 32452
rect 5236 32396 6412 32452
rect 6468 32396 9436 32452
rect 9492 32396 9502 32452
rect 25554 32396 25564 32452
rect 25620 32396 27916 32452
rect 27972 32396 27982 32452
rect 37874 32396 37884 32452
rect 37940 32396 39340 32452
rect 39396 32396 39406 32452
rect 43922 32396 43932 32452
rect 43988 32396 49084 32452
rect 49140 32396 49150 32452
rect 30818 32284 30828 32340
rect 30884 32284 35644 32340
rect 35700 32284 35710 32340
rect 45042 32284 45052 32340
rect 45108 32284 48860 32340
rect 48916 32284 48926 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 28578 32060 28588 32116
rect 28644 32060 34916 32116
rect 34860 32004 34916 32060
rect 38612 32060 42028 32116
rect 42084 32060 42094 32116
rect 38612 32004 38668 32060
rect 13468 31948 13972 32004
rect 14130 31948 14140 32004
rect 14196 31948 15148 32004
rect 15204 31948 15214 32004
rect 31154 31948 31164 32004
rect 31220 31948 34636 32004
rect 34692 31948 34702 32004
rect 34860 31948 38668 32004
rect 39218 31948 39228 32004
rect 39284 31948 40124 32004
rect 40180 31948 40190 32004
rect 13468 31892 13524 31948
rect 13916 31892 13972 31948
rect 2482 31836 2492 31892
rect 2548 31836 5852 31892
rect 5908 31836 5918 31892
rect 6290 31836 6300 31892
rect 6356 31836 7532 31892
rect 7588 31836 10892 31892
rect 10948 31836 13524 31892
rect 13682 31836 13692 31892
rect 13748 31836 13758 31892
rect 13916 31836 43820 31892
rect 43876 31836 43886 31892
rect 50530 31836 50540 31892
rect 50596 31836 52444 31892
rect 52500 31836 52510 31892
rect 13692 31780 13748 31836
rect 13692 31724 21868 31780
rect 21924 31724 23548 31780
rect 23604 31724 23614 31780
rect 29474 31724 29484 31780
rect 29540 31724 31724 31780
rect 31780 31724 32284 31780
rect 32340 31724 32350 31780
rect 39218 31724 39228 31780
rect 39284 31724 39900 31780
rect 39956 31724 43372 31780
rect 43428 31724 43438 31780
rect 4722 31612 4732 31668
rect 4788 31612 5292 31668
rect 5348 31612 5358 31668
rect 16146 31612 16156 31668
rect 16212 31612 16604 31668
rect 16660 31612 16670 31668
rect 19170 31612 19180 31668
rect 19236 31612 21532 31668
rect 21588 31612 23660 31668
rect 23716 31612 23726 31668
rect 24994 31612 25004 31668
rect 25060 31612 39396 31668
rect 45266 31612 45276 31668
rect 45332 31612 46396 31668
rect 46452 31612 46462 31668
rect 5058 31500 5068 31556
rect 5124 31500 6748 31556
rect 6804 31500 8204 31556
rect 8260 31500 15932 31556
rect 15988 31500 15998 31556
rect 26002 31500 26012 31556
rect 26068 31500 26460 31556
rect 26516 31500 26526 31556
rect 28130 31500 28140 31556
rect 28196 31500 28588 31556
rect 28644 31500 29260 31556
rect 29316 31500 29708 31556
rect 29764 31500 35532 31556
rect 35588 31500 35598 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 26460 31220 26516 31500
rect 39340 31444 39396 31612
rect 39554 31500 39564 31556
rect 39620 31500 42812 31556
rect 42868 31500 42878 31556
rect 49858 31500 49868 31556
rect 49924 31500 50428 31556
rect 50484 31500 51100 31556
rect 51156 31500 51166 31556
rect 30482 31388 30492 31444
rect 30548 31388 31612 31444
rect 31668 31388 31678 31444
rect 39340 31388 43372 31444
rect 43428 31388 43438 31444
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 26674 31276 26684 31332
rect 26740 31276 27020 31332
rect 27076 31276 27468 31332
rect 27524 31276 27534 31332
rect 29586 31276 29596 31332
rect 29652 31276 38668 31332
rect 38612 31220 38668 31276
rect 16370 31164 16380 31220
rect 16436 31164 17724 31220
rect 17780 31164 21084 31220
rect 21140 31164 22764 31220
rect 22820 31164 22830 31220
rect 26460 31164 29932 31220
rect 29988 31164 29998 31220
rect 38612 31164 40348 31220
rect 40404 31164 40414 31220
rect 43810 31164 43820 31220
rect 43876 31164 44828 31220
rect 44884 31164 44894 31220
rect 20402 31052 20412 31108
rect 20468 31052 21644 31108
rect 21700 31052 21710 31108
rect 22194 31052 22204 31108
rect 22260 31052 22988 31108
rect 23044 31052 23054 31108
rect 25442 31052 25452 31108
rect 25508 31052 34300 31108
rect 34356 31052 35308 31108
rect 35364 31052 35374 31108
rect 35522 31052 35532 31108
rect 35588 31052 42140 31108
rect 42196 31052 42206 31108
rect 44370 31052 44380 31108
rect 44436 31052 45052 31108
rect 45108 31052 45118 31108
rect 5618 30940 5628 30996
rect 5684 30940 6300 30996
rect 6356 30940 6366 30996
rect 9874 30940 9884 30996
rect 9940 30940 10220 30996
rect 10276 30940 10286 30996
rect 16482 30940 16492 30996
rect 16548 30940 16716 30996
rect 16772 30940 16782 30996
rect 21522 30940 21532 30996
rect 21588 30940 22316 30996
rect 22372 30940 22382 30996
rect 26450 30940 26460 30996
rect 26516 30940 27692 30996
rect 27748 30940 27758 30996
rect 28130 30940 28140 30996
rect 28196 30940 31276 30996
rect 31332 30940 31342 30996
rect 28140 30884 28196 30940
rect 35308 30884 35364 31052
rect 16370 30828 16380 30884
rect 16436 30828 16940 30884
rect 16996 30828 17006 30884
rect 18274 30828 18284 30884
rect 18340 30828 22540 30884
rect 22596 30828 23884 30884
rect 23940 30828 23950 30884
rect 27570 30828 27580 30884
rect 27636 30828 28196 30884
rect 30818 30828 30828 30884
rect 30884 30828 33068 30884
rect 33124 30828 33134 30884
rect 35308 30828 39004 30884
rect 39060 30828 39070 30884
rect 48962 30828 48972 30884
rect 49028 30828 49980 30884
rect 50036 30828 50046 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 4610 30268 4620 30324
rect 4676 30268 5740 30324
rect 5796 30268 5806 30324
rect 6748 30268 7196 30324
rect 7252 30268 8316 30324
rect 8372 30268 8382 30324
rect 17938 30268 17948 30324
rect 18004 30268 19404 30324
rect 19460 30268 26012 30324
rect 26068 30268 26078 30324
rect 42130 30268 42140 30324
rect 42196 30268 43372 30324
rect 43428 30268 43438 30324
rect 49634 30268 49644 30324
rect 49700 30268 52892 30324
rect 52948 30268 52958 30324
rect 6748 30100 6804 30268
rect 6962 30156 6972 30212
rect 7028 30156 7756 30212
rect 7812 30156 8652 30212
rect 8708 30156 8718 30212
rect 15092 30156 18172 30212
rect 18228 30156 18238 30212
rect 21746 30156 21756 30212
rect 21812 30156 22316 30212
rect 22372 30156 22382 30212
rect 24098 30156 24108 30212
rect 24164 30156 25004 30212
rect 25060 30156 28700 30212
rect 28756 30156 29148 30212
rect 29204 30156 29214 30212
rect 31378 30156 31388 30212
rect 31444 30156 31612 30212
rect 31668 30156 34188 30212
rect 34244 30156 34254 30212
rect 42578 30156 42588 30212
rect 42644 30156 43148 30212
rect 43204 30156 43214 30212
rect 15092 30100 15148 30156
rect 54200 30100 55000 30128
rect 2482 30044 2492 30100
rect 2548 30044 6300 30100
rect 6356 30044 6366 30100
rect 6738 30044 6748 30100
rect 6804 30044 6814 30100
rect 8418 30044 8428 30100
rect 8484 30044 15148 30100
rect 15810 30044 15820 30100
rect 15876 30044 17276 30100
rect 17332 30044 17342 30100
rect 22530 30044 22540 30100
rect 22596 30044 23100 30100
rect 23156 30044 25452 30100
rect 25508 30044 25518 30100
rect 29698 30044 29708 30100
rect 29764 30044 30268 30100
rect 30324 30044 30334 30100
rect 53218 30044 53228 30100
rect 53284 30044 55000 30100
rect 54200 30016 55000 30044
rect 26338 29932 26348 29988
rect 26404 29932 27020 29988
rect 27076 29932 31276 29988
rect 31332 29932 31948 29988
rect 32004 29932 32508 29988
rect 32564 29932 32574 29988
rect 34850 29932 34860 29988
rect 34916 29932 34926 29988
rect 35634 29932 35644 29988
rect 35700 29932 36876 29988
rect 36932 29932 39452 29988
rect 39508 29932 40572 29988
rect 40628 29932 41356 29988
rect 41412 29932 41422 29988
rect 43138 29932 43148 29988
rect 43204 29932 45164 29988
rect 45220 29932 45724 29988
rect 45780 29932 48300 29988
rect 48356 29932 48366 29988
rect 34860 29876 34916 29932
rect 21074 29820 21084 29876
rect 21140 29820 21980 29876
rect 22036 29820 33740 29876
rect 33796 29820 35868 29876
rect 35924 29820 35934 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 6860 29708 7084 29764
rect 7140 29708 7150 29764
rect 30594 29708 30604 29764
rect 30660 29708 31724 29764
rect 31780 29708 34076 29764
rect 34132 29708 34142 29764
rect 39302 29708 39340 29764
rect 39396 29708 39406 29764
rect 6860 29652 6916 29708
rect 6850 29596 6860 29652
rect 6916 29596 6926 29652
rect 12898 29596 12908 29652
rect 12964 29596 13692 29652
rect 13748 29596 13758 29652
rect 17266 29596 17276 29652
rect 17332 29596 22652 29652
rect 22708 29596 22718 29652
rect 27906 29596 27916 29652
rect 27972 29596 29596 29652
rect 29652 29596 29662 29652
rect 35074 29596 35084 29652
rect 35140 29596 35980 29652
rect 36036 29596 39228 29652
rect 39284 29596 39294 29652
rect 42018 29596 42028 29652
rect 42084 29596 43820 29652
rect 43876 29596 45500 29652
rect 45556 29596 45566 29652
rect 23762 29484 23772 29540
rect 23828 29484 26908 29540
rect 26964 29484 26974 29540
rect 33506 29484 33516 29540
rect 33572 29484 34972 29540
rect 35028 29484 35532 29540
rect 35588 29484 38668 29540
rect 48178 29484 48188 29540
rect 48244 29484 51212 29540
rect 51268 29484 51278 29540
rect 6402 29372 6412 29428
rect 6468 29372 6748 29428
rect 6804 29372 6814 29428
rect 8866 29372 8876 29428
rect 8932 29372 9548 29428
rect 9604 29372 10780 29428
rect 10836 29372 10846 29428
rect 26852 29372 30828 29428
rect 30884 29372 32172 29428
rect 32228 29372 34300 29428
rect 34356 29372 37100 29428
rect 37156 29372 37166 29428
rect 26852 29316 26908 29372
rect 8978 29260 8988 29316
rect 9044 29260 9884 29316
rect 9940 29260 10444 29316
rect 10500 29260 10510 29316
rect 10882 29260 10892 29316
rect 10948 29260 12684 29316
rect 12740 29260 12750 29316
rect 13010 29260 13020 29316
rect 13076 29260 14140 29316
rect 14196 29260 14206 29316
rect 15474 29260 15484 29316
rect 15540 29260 16828 29316
rect 16884 29260 17724 29316
rect 17780 29260 17790 29316
rect 18834 29260 18844 29316
rect 18900 29260 22876 29316
rect 22932 29260 26908 29316
rect 28018 29260 28028 29316
rect 28084 29260 28812 29316
rect 28868 29260 28878 29316
rect 38612 29092 38668 29484
rect 40450 29372 40460 29428
rect 40516 29372 41132 29428
rect 41188 29372 41198 29428
rect 47058 29372 47068 29428
rect 47124 29372 47964 29428
rect 48020 29372 48030 29428
rect 49970 29372 49980 29428
rect 50036 29372 51884 29428
rect 51940 29372 52444 29428
rect 52500 29372 53116 29428
rect 53172 29372 53182 29428
rect 39890 29260 39900 29316
rect 39956 29260 42700 29316
rect 42756 29260 42766 29316
rect 12114 29036 12124 29092
rect 12180 29036 12190 29092
rect 16258 29036 16268 29092
rect 16324 29036 17724 29092
rect 17780 29036 17790 29092
rect 38612 29036 40012 29092
rect 40068 29036 40078 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 12124 28980 12180 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 12124 28924 12796 28980
rect 12852 28924 19628 28980
rect 19684 28924 19694 28980
rect 12898 28812 12908 28868
rect 12964 28812 13356 28868
rect 13412 28812 17668 28868
rect 27122 28812 27132 28868
rect 27188 28812 28140 28868
rect 28196 28812 42588 28868
rect 42644 28812 42654 28868
rect 43474 28812 43484 28868
rect 43540 28812 47068 28868
rect 47124 28812 47964 28868
rect 48020 28812 49084 28868
rect 49140 28812 49150 28868
rect 9650 28700 9660 28756
rect 9716 28700 10220 28756
rect 10276 28700 11340 28756
rect 11396 28700 11900 28756
rect 11956 28700 11966 28756
rect 13458 28700 13468 28756
rect 13524 28700 16492 28756
rect 16548 28700 16558 28756
rect 17612 28644 17668 28812
rect 18162 28700 18172 28756
rect 18228 28700 18732 28756
rect 18788 28700 18798 28756
rect 20066 28700 20076 28756
rect 20132 28700 20748 28756
rect 20804 28700 20814 28756
rect 22642 28700 22652 28756
rect 22708 28700 23212 28756
rect 23268 28700 23278 28756
rect 31378 28700 31388 28756
rect 31444 28700 33628 28756
rect 33684 28700 34972 28756
rect 35028 28700 35038 28756
rect 36642 28700 36652 28756
rect 36708 28700 37324 28756
rect 37380 28700 37390 28756
rect 48290 28700 48300 28756
rect 48356 28700 48972 28756
rect 49028 28700 49038 28756
rect 5730 28588 5740 28644
rect 5796 28588 8428 28644
rect 8484 28588 8494 28644
rect 12460 28588 16268 28644
rect 16324 28588 16334 28644
rect 17602 28588 17612 28644
rect 17668 28588 17678 28644
rect 27570 28588 27580 28644
rect 27636 28588 28028 28644
rect 28084 28588 28094 28644
rect 36530 28588 36540 28644
rect 36596 28588 37212 28644
rect 37268 28588 37278 28644
rect 37986 28588 37996 28644
rect 38052 28588 38780 28644
rect 38836 28588 38846 28644
rect 38994 28588 39004 28644
rect 39060 28588 40572 28644
rect 40628 28588 41356 28644
rect 41412 28588 41422 28644
rect 48300 28588 49084 28644
rect 49140 28588 49150 28644
rect 12460 28532 12516 28588
rect 6402 28476 6412 28532
rect 6468 28476 7196 28532
rect 7252 28476 7262 28532
rect 10658 28476 10668 28532
rect 10724 28476 11452 28532
rect 11508 28476 12460 28532
rect 12516 28476 12526 28532
rect 21858 28476 21868 28532
rect 21924 28476 22540 28532
rect 22596 28476 25676 28532
rect 25732 28476 25742 28532
rect 28578 28476 28588 28532
rect 28644 28476 30044 28532
rect 30100 28476 31724 28532
rect 31780 28476 32732 28532
rect 32788 28476 32798 28532
rect 40236 28420 40292 28588
rect 40786 28476 40796 28532
rect 40852 28476 41804 28532
rect 41860 28476 42700 28532
rect 42756 28476 42766 28532
rect 46498 28476 46508 28532
rect 46564 28476 48076 28532
rect 48132 28476 48142 28532
rect 48300 28420 48356 28588
rect 23202 28364 23212 28420
rect 23268 28364 26012 28420
rect 26068 28364 26460 28420
rect 26516 28364 26526 28420
rect 27906 28364 27916 28420
rect 27972 28364 30492 28420
rect 30548 28364 30828 28420
rect 30884 28364 30894 28420
rect 40226 28364 40236 28420
rect 40292 28364 40302 28420
rect 41010 28364 41020 28420
rect 41076 28364 48356 28420
rect 24658 28252 24668 28308
rect 24724 28252 33516 28308
rect 33572 28252 33582 28308
rect 38994 28252 39004 28308
rect 39060 28252 39452 28308
rect 39508 28252 44716 28308
rect 44772 28252 44782 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 20962 28140 20972 28196
rect 21028 28140 26796 28196
rect 26852 28140 27916 28196
rect 27972 28140 27982 28196
rect 28242 28140 28252 28196
rect 28308 28140 29708 28196
rect 29764 28140 29774 28196
rect 34514 28140 34524 28196
rect 34580 28140 35196 28196
rect 35252 28140 35532 28196
rect 35588 28140 35598 28196
rect 5282 28028 5292 28084
rect 5348 28028 5964 28084
rect 6020 28028 6030 28084
rect 6178 28028 6188 28084
rect 6244 28028 6636 28084
rect 6692 28028 6702 28084
rect 7522 28028 7532 28084
rect 7588 28028 9324 28084
rect 9380 28028 9390 28084
rect 19618 28028 19628 28084
rect 19684 28028 20300 28084
rect 20356 28028 20636 28084
rect 20692 28028 20702 28084
rect 22642 28028 22652 28084
rect 22708 28028 34972 28084
rect 35028 28028 35980 28084
rect 36036 28028 36046 28084
rect 39106 28028 39116 28084
rect 39172 28028 39564 28084
rect 39620 28028 39630 28084
rect 40002 28028 40012 28084
rect 40068 28028 40236 28084
rect 40292 28028 41020 28084
rect 41076 28028 41086 28084
rect 6066 27916 6076 27972
rect 6132 27916 7756 27972
rect 7812 27916 7822 27972
rect 24098 27916 24108 27972
rect 24164 27916 24668 27972
rect 24724 27916 24734 27972
rect 30370 27916 30380 27972
rect 30436 27916 31276 27972
rect 31332 27916 31342 27972
rect 4946 27804 4956 27860
rect 5012 27804 8540 27860
rect 8596 27804 19068 27860
rect 19124 27804 19134 27860
rect 22418 27804 22428 27860
rect 22484 27804 24220 27860
rect 24276 27804 24286 27860
rect 33954 27804 33964 27860
rect 34020 27804 34748 27860
rect 34804 27804 34814 27860
rect 35634 27804 35644 27860
rect 35700 27804 44268 27860
rect 44324 27804 45052 27860
rect 45108 27804 45118 27860
rect 48188 27804 48636 27860
rect 48692 27804 48702 27860
rect 48188 27748 48244 27804
rect 2482 27692 2492 27748
rect 2548 27692 6860 27748
rect 6916 27692 6926 27748
rect 13906 27692 13916 27748
rect 13972 27692 26908 27748
rect 26964 27692 27244 27748
rect 27300 27692 27310 27748
rect 38098 27692 38108 27748
rect 38164 27692 38556 27748
rect 38612 27692 39340 27748
rect 39396 27692 39406 27748
rect 41458 27692 41468 27748
rect 41524 27692 44604 27748
rect 44660 27692 48244 27748
rect 48402 27692 48412 27748
rect 48468 27692 49980 27748
rect 50036 27692 50046 27748
rect 6514 27580 6524 27636
rect 6580 27580 8316 27636
rect 8372 27580 8382 27636
rect 21970 27580 21980 27636
rect 22036 27580 23324 27636
rect 23380 27580 23390 27636
rect 35970 27468 35980 27524
rect 36036 27468 40236 27524
rect 40292 27468 40302 27524
rect 45602 27468 45612 27524
rect 45668 27468 45948 27524
rect 46004 27468 47628 27524
rect 47684 27468 47694 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 54200 27412 55000 27440
rect 32722 27356 32732 27412
rect 32788 27356 34188 27412
rect 34244 27356 34254 27412
rect 39330 27356 39340 27412
rect 39396 27356 39676 27412
rect 39732 27356 40684 27412
rect 40740 27356 40750 27412
rect 53330 27356 53340 27412
rect 53396 27356 55000 27412
rect 54200 27328 55000 27356
rect 6626 27244 6636 27300
rect 6692 27244 7308 27300
rect 7364 27244 7374 27300
rect 10994 27244 11004 27300
rect 11060 27244 11070 27300
rect 25666 27244 25676 27300
rect 25732 27244 27580 27300
rect 27636 27244 27646 27300
rect 31042 27244 31052 27300
rect 31108 27244 31836 27300
rect 31892 27244 37100 27300
rect 37156 27244 37166 27300
rect 43698 27244 43708 27300
rect 43764 27244 45052 27300
rect 45108 27244 45118 27300
rect 47058 27244 47068 27300
rect 47124 27244 47516 27300
rect 47572 27244 47582 27300
rect 51650 27244 51660 27300
rect 51716 27244 52444 27300
rect 52500 27244 52510 27300
rect 5282 27132 5292 27188
rect 5348 27132 6524 27188
rect 6580 27132 6590 27188
rect 11004 26964 11060 27244
rect 23202 27132 23212 27188
rect 23268 27132 23884 27188
rect 23940 27132 23950 27188
rect 30678 27132 30716 27188
rect 30772 27132 32284 27188
rect 32340 27132 36092 27188
rect 36148 27132 46508 27188
rect 46564 27132 46574 27188
rect 22306 27020 22316 27076
rect 22372 27020 22596 27076
rect 31938 27020 31948 27076
rect 32004 27020 34524 27076
rect 34580 27020 35644 27076
rect 35700 27020 35710 27076
rect 35858 27020 35868 27076
rect 35924 27020 36316 27076
rect 36372 27020 36382 27076
rect 37202 27020 37212 27076
rect 37268 27020 39228 27076
rect 39284 27020 39294 27076
rect 40674 27020 40684 27076
rect 40740 27020 41468 27076
rect 41524 27020 41534 27076
rect 22540 26964 22596 27020
rect 11004 26908 11284 26964
rect 12898 26908 12908 26964
rect 12964 26908 14252 26964
rect 14308 26908 14318 26964
rect 21634 26908 21644 26964
rect 21700 26908 22204 26964
rect 22260 26908 22270 26964
rect 22530 26908 22540 26964
rect 22596 26908 22606 26964
rect 29026 26908 29036 26964
rect 29092 26908 30604 26964
rect 30660 26908 30670 26964
rect 31602 26908 31612 26964
rect 31668 26908 34412 26964
rect 34468 26908 34860 26964
rect 34916 26908 34926 26964
rect 37650 26908 37660 26964
rect 37716 26908 38444 26964
rect 38500 26908 39116 26964
rect 39172 26908 40012 26964
rect 40068 26908 40078 26964
rect 40338 26908 40348 26964
rect 40404 26908 41020 26964
rect 41076 26908 44604 26964
rect 44660 26908 44670 26964
rect 11228 26852 11284 26908
rect 10994 26796 11004 26852
rect 11060 26796 11284 26852
rect 27570 26796 27580 26852
rect 27636 26796 29148 26852
rect 29204 26796 37100 26852
rect 37156 26796 37884 26852
rect 37940 26796 37950 26852
rect 44370 26796 44380 26852
rect 44436 26796 44828 26852
rect 44884 26796 44894 26852
rect 12002 26684 12012 26740
rect 12068 26684 12078 26740
rect 27682 26684 27692 26740
rect 27748 26684 28140 26740
rect 28196 26684 28206 26740
rect 5842 26460 5852 26516
rect 5908 26460 6636 26516
rect 6692 26460 6702 26516
rect 12012 26404 12068 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 20626 26572 20636 26628
rect 20692 26572 28924 26628
rect 28980 26572 28990 26628
rect 39974 26572 40012 26628
rect 40068 26572 40078 26628
rect 27570 26460 27580 26516
rect 27636 26460 28028 26516
rect 28084 26460 28094 26516
rect 38612 26460 39900 26516
rect 39956 26460 39966 26516
rect 12012 26348 15260 26404
rect 15316 26348 15326 26404
rect 30258 26348 30268 26404
rect 30324 26348 30334 26404
rect 6066 26236 6076 26292
rect 6132 26236 6524 26292
rect 6580 26236 6972 26292
rect 7028 26236 7038 26292
rect 11218 26236 11228 26292
rect 11284 26236 12348 26292
rect 12404 26236 12414 26292
rect 12572 26180 12628 26348
rect 30268 26292 30324 26348
rect 24434 26236 24444 26292
rect 24500 26236 25900 26292
rect 25956 26236 25966 26292
rect 30268 26236 30828 26292
rect 30884 26236 30894 26292
rect 11778 26124 11788 26180
rect 11844 26124 12628 26180
rect 18274 26124 18284 26180
rect 18340 26124 18844 26180
rect 18900 26124 28588 26180
rect 28644 26124 28654 26180
rect 29810 26124 29820 26180
rect 29876 26124 30268 26180
rect 30324 26124 31276 26180
rect 31332 26124 31342 26180
rect 38612 26068 38668 26460
rect 45154 26348 45164 26404
rect 45220 26348 49868 26404
rect 49924 26348 52892 26404
rect 52948 26348 52958 26404
rect 39890 26124 39900 26180
rect 39956 26124 43036 26180
rect 43092 26124 43102 26180
rect 43810 26124 43820 26180
rect 43876 26124 44268 26180
rect 44324 26124 45388 26180
rect 45444 26124 45454 26180
rect 10994 26012 11004 26068
rect 11060 26012 11900 26068
rect 11956 26012 11966 26068
rect 38322 26012 38332 26068
rect 38388 26012 38668 26068
rect 49858 26012 49868 26068
rect 49924 26012 51660 26068
rect 51716 26012 51726 26068
rect 11554 25900 11564 25956
rect 11620 25900 12348 25956
rect 12404 25900 12414 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 18386 25676 18396 25732
rect 18452 25676 19628 25732
rect 19684 25676 19694 25732
rect 21634 25676 21644 25732
rect 21700 25676 22316 25732
rect 22372 25676 22382 25732
rect 27122 25676 27132 25732
rect 27188 25676 31164 25732
rect 31220 25676 32172 25732
rect 32228 25676 34860 25732
rect 34916 25676 34926 25732
rect 6066 25564 6076 25620
rect 6132 25564 9324 25620
rect 9380 25564 9660 25620
rect 9716 25564 9726 25620
rect 31714 25564 31724 25620
rect 31780 25564 31948 25620
rect 32004 25564 32014 25620
rect 35074 25564 35084 25620
rect 35140 25564 36428 25620
rect 36484 25564 38332 25620
rect 38388 25564 38398 25620
rect 5394 25452 5404 25508
rect 5460 25452 5628 25508
rect 5684 25452 9436 25508
rect 9492 25452 17948 25508
rect 18004 25452 18014 25508
rect 18610 25452 18620 25508
rect 18676 25452 19516 25508
rect 19572 25452 19582 25508
rect 25890 25452 25900 25508
rect 25956 25452 26908 25508
rect 27906 25452 27916 25508
rect 27972 25452 29372 25508
rect 29428 25452 30492 25508
rect 30548 25452 43708 25508
rect 43764 25452 44268 25508
rect 44324 25452 44334 25508
rect 49858 25452 49868 25508
rect 49924 25452 51100 25508
rect 51156 25452 51166 25508
rect 9538 25340 9548 25396
rect 9604 25340 10332 25396
rect 10388 25340 10398 25396
rect 10658 25340 10668 25396
rect 10724 25340 11340 25396
rect 11396 25340 11406 25396
rect 2930 25228 2940 25284
rect 2996 25228 5964 25284
rect 6020 25228 6030 25284
rect 11340 25172 11396 25340
rect 18386 25228 18396 25284
rect 18452 25228 19068 25284
rect 19124 25228 19134 25284
rect 25554 25228 25564 25284
rect 25620 25228 26572 25284
rect 26628 25228 26638 25284
rect 26852 25228 26908 25452
rect 28130 25340 28140 25396
rect 28196 25340 29932 25396
rect 29988 25340 38668 25396
rect 49522 25340 49532 25396
rect 49588 25340 50204 25396
rect 50260 25340 50270 25396
rect 38612 25284 38668 25340
rect 26964 25228 28476 25284
rect 28532 25228 28542 25284
rect 31266 25228 31276 25284
rect 31332 25228 33628 25284
rect 33684 25228 34748 25284
rect 34804 25228 35532 25284
rect 35588 25228 35598 25284
rect 38612 25228 40796 25284
rect 40852 25228 40862 25284
rect 43362 25228 43372 25284
rect 43428 25228 44268 25284
rect 44324 25228 44334 25284
rect 46946 25228 46956 25284
rect 47012 25228 50540 25284
rect 50596 25228 50606 25284
rect 11330 25116 11340 25172
rect 11396 25116 11406 25172
rect 26450 25116 26460 25172
rect 26516 25116 27132 25172
rect 27188 25116 27198 25172
rect 34962 25116 34972 25172
rect 35028 25116 36316 25172
rect 36372 25116 39676 25172
rect 39732 25116 39742 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 50988 24948 51044 25452
rect 51314 25116 51324 25172
rect 51380 25116 51390 25172
rect 13122 24892 13132 24948
rect 13188 24892 14700 24948
rect 14756 24892 14766 24948
rect 18946 24892 18956 24948
rect 19012 24892 20188 24948
rect 20244 24892 21308 24948
rect 21364 24892 21374 24948
rect 28578 24892 28588 24948
rect 28644 24892 30268 24948
rect 30324 24892 30716 24948
rect 30772 24892 30782 24948
rect 31042 24892 31052 24948
rect 31108 24892 41244 24948
rect 41300 24892 41310 24948
rect 50754 24892 50764 24948
rect 50820 24892 51044 24948
rect 51324 24836 51380 25116
rect 11666 24780 11676 24836
rect 11732 24780 13580 24836
rect 13636 24780 16828 24836
rect 16884 24780 16894 24836
rect 19058 24780 19068 24836
rect 19124 24780 22540 24836
rect 22596 24780 25564 24836
rect 25620 24780 25630 24836
rect 26114 24780 26124 24836
rect 26180 24780 28364 24836
rect 28420 24780 28430 24836
rect 28914 24780 28924 24836
rect 28980 24780 29708 24836
rect 29764 24780 30604 24836
rect 30660 24780 32060 24836
rect 32116 24780 32396 24836
rect 32452 24780 32462 24836
rect 37986 24780 37996 24836
rect 38052 24780 39060 24836
rect 43810 24780 43820 24836
rect 43876 24780 46284 24836
rect 46340 24780 46350 24836
rect 50866 24780 50876 24836
rect 50932 24780 51380 24836
rect 39004 24724 39060 24780
rect 54200 24724 55000 24752
rect 4610 24668 4620 24724
rect 4676 24668 5404 24724
rect 5460 24668 5470 24724
rect 12674 24668 12684 24724
rect 12740 24668 13468 24724
rect 13524 24668 13534 24724
rect 16706 24668 16716 24724
rect 16772 24668 18284 24724
rect 18340 24668 18350 24724
rect 22978 24668 22988 24724
rect 23044 24668 23660 24724
rect 23716 24668 23726 24724
rect 28140 24668 29036 24724
rect 29092 24668 29102 24724
rect 35522 24668 35532 24724
rect 35588 24668 38780 24724
rect 38836 24668 38846 24724
rect 38994 24668 39004 24724
rect 39060 24668 40348 24724
rect 40404 24668 41244 24724
rect 41300 24668 41310 24724
rect 48738 24668 48748 24724
rect 48804 24668 49420 24724
rect 49476 24668 49868 24724
rect 49924 24668 49934 24724
rect 50306 24668 50316 24724
rect 50372 24668 51660 24724
rect 51716 24668 51726 24724
rect 53218 24668 53228 24724
rect 53284 24668 55000 24724
rect 28140 24612 28196 24668
rect 49868 24612 49924 24668
rect 54200 24640 55000 24668
rect 11666 24556 11676 24612
rect 11732 24556 12796 24612
rect 12852 24556 12862 24612
rect 26898 24556 26908 24612
rect 26964 24556 27468 24612
rect 27524 24556 28140 24612
rect 28196 24556 28206 24612
rect 32610 24556 32620 24612
rect 32676 24556 34636 24612
rect 34692 24556 34702 24612
rect 37986 24556 37996 24612
rect 38052 24556 39340 24612
rect 39396 24556 39406 24612
rect 48178 24556 48188 24612
rect 48244 24556 48860 24612
rect 48916 24556 48926 24612
rect 49868 24556 50204 24612
rect 50260 24556 50270 24612
rect 44034 24444 44044 24500
rect 44100 24444 44828 24500
rect 44884 24444 44894 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 24770 23996 24780 24052
rect 24836 23996 26236 24052
rect 26292 23996 26302 24052
rect 34962 23996 34972 24052
rect 35028 23996 37268 24052
rect 37212 23940 37268 23996
rect 34402 23884 34412 23940
rect 34468 23884 35644 23940
rect 35700 23884 35710 23940
rect 37202 23884 37212 23940
rect 37268 23884 38556 23940
rect 38612 23884 38622 23940
rect 44258 23884 44268 23940
rect 44324 23884 45052 23940
rect 45108 23884 45118 23940
rect 49858 23884 49868 23940
rect 49924 23884 50428 23940
rect 50484 23884 50494 23940
rect 35970 23772 35980 23828
rect 36036 23772 36876 23828
rect 36932 23772 36942 23828
rect 46274 23772 46284 23828
rect 46340 23772 46732 23828
rect 46788 23772 52108 23828
rect 52164 23772 52174 23828
rect 2706 23660 2716 23716
rect 2772 23660 3388 23716
rect 3444 23660 3454 23716
rect 5954 23660 5964 23716
rect 6020 23660 6636 23716
rect 6692 23660 6702 23716
rect 37090 23660 37100 23716
rect 37156 23660 38332 23716
rect 38388 23660 38398 23716
rect 45714 23660 45724 23716
rect 45780 23660 47404 23716
rect 47460 23660 47470 23716
rect 49298 23660 49308 23716
rect 49364 23660 49756 23716
rect 49812 23660 52892 23716
rect 52948 23660 52958 23716
rect 10434 23548 10444 23604
rect 10500 23548 11228 23604
rect 11284 23548 11294 23604
rect 40002 23548 40012 23604
rect 40068 23548 40908 23604
rect 40964 23548 40974 23604
rect 43810 23548 43820 23604
rect 43876 23548 44268 23604
rect 44324 23548 44334 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 7186 23436 7196 23492
rect 7252 23436 8092 23492
rect 8148 23436 10220 23492
rect 10276 23436 10286 23492
rect 11330 23436 11340 23492
rect 11396 23436 13356 23492
rect 13412 23436 18788 23492
rect 38098 23436 38108 23492
rect 38164 23436 39788 23492
rect 39844 23436 39854 23492
rect 10098 23324 10108 23380
rect 10164 23324 11452 23380
rect 11508 23324 12908 23380
rect 12964 23324 18508 23380
rect 18564 23324 18574 23380
rect 18732 23268 18788 23436
rect 44930 23324 44940 23380
rect 44996 23324 45388 23380
rect 45444 23324 48412 23380
rect 48468 23324 49196 23380
rect 49252 23324 50428 23380
rect 11554 23212 11564 23268
rect 11620 23212 12684 23268
rect 12740 23212 12750 23268
rect 18274 23212 18284 23268
rect 18340 23212 20524 23268
rect 20580 23212 20590 23268
rect 39442 23212 39452 23268
rect 39508 23212 41356 23268
rect 41412 23212 41422 23268
rect 41794 23212 41804 23268
rect 41860 23212 42700 23268
rect 42756 23212 43036 23268
rect 43092 23212 43102 23268
rect 50372 23156 50428 23324
rect 13010 23100 13020 23156
rect 13076 23100 14364 23156
rect 14420 23100 14430 23156
rect 14914 23100 14924 23156
rect 14980 23100 19516 23156
rect 19572 23100 19582 23156
rect 20402 23100 20412 23156
rect 20468 23100 21196 23156
rect 21252 23100 24780 23156
rect 24836 23100 24846 23156
rect 36754 23100 36764 23156
rect 36820 23100 48748 23156
rect 48804 23100 48814 23156
rect 50372 23100 50876 23156
rect 50932 23100 53116 23156
rect 53172 23100 53182 23156
rect 7522 22988 7532 23044
rect 7588 22988 13244 23044
rect 13300 22988 13310 23044
rect 26002 22988 26012 23044
rect 26068 22988 27356 23044
rect 27412 22988 28588 23044
rect 28644 22988 28654 23044
rect 42130 22988 42140 23044
rect 42196 22988 43036 23044
rect 43092 22988 43484 23044
rect 43540 22988 43550 23044
rect 11554 22876 11564 22932
rect 11620 22876 14028 22932
rect 14084 22876 14094 22932
rect 37202 22876 37212 22932
rect 37268 22876 39116 22932
rect 39172 22876 39182 22932
rect 39666 22876 39676 22932
rect 39732 22876 41804 22932
rect 41860 22876 41870 22932
rect 42578 22876 42588 22932
rect 42644 22876 44044 22932
rect 44100 22876 45388 22932
rect 45444 22876 45454 22932
rect 42588 22820 42644 22876
rect 41234 22764 41244 22820
rect 41300 22764 42644 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 29250 22652 29260 22708
rect 29316 22652 31500 22708
rect 31556 22652 31566 22708
rect 8306 22540 8316 22596
rect 8372 22540 10668 22596
rect 10724 22540 10734 22596
rect 14354 22540 14364 22596
rect 14420 22540 15372 22596
rect 15428 22540 15932 22596
rect 15988 22540 15998 22596
rect 13010 22428 13020 22484
rect 13076 22428 13692 22484
rect 13748 22428 13758 22484
rect 15092 22428 29148 22484
rect 29204 22428 29214 22484
rect 31154 22428 31164 22484
rect 31220 22428 37100 22484
rect 37156 22428 37166 22484
rect 47954 22428 47964 22484
rect 48020 22428 49196 22484
rect 49252 22428 49262 22484
rect 15092 22372 15148 22428
rect 5170 22316 5180 22372
rect 5236 22316 7084 22372
rect 7140 22316 7150 22372
rect 7634 22316 7644 22372
rect 7700 22316 8316 22372
rect 8372 22316 8988 22372
rect 9044 22316 9054 22372
rect 10770 22316 10780 22372
rect 10836 22316 11900 22372
rect 11956 22316 13132 22372
rect 13188 22316 13198 22372
rect 13906 22316 13916 22372
rect 13972 22316 14812 22372
rect 14868 22316 15148 22372
rect 23650 22316 23660 22372
rect 23716 22316 24332 22372
rect 24388 22316 26012 22372
rect 26068 22316 26078 22372
rect 5852 22260 5908 22316
rect 5842 22204 5852 22260
rect 5908 22204 5918 22260
rect 7746 22204 7756 22260
rect 7812 22204 7980 22260
rect 8036 22204 8764 22260
rect 8820 22204 8830 22260
rect 9314 22204 9324 22260
rect 9380 22204 9996 22260
rect 10052 22204 13468 22260
rect 13524 22204 13534 22260
rect 18946 22204 18956 22260
rect 19012 22204 20636 22260
rect 20692 22204 20702 22260
rect 24994 22204 25004 22260
rect 25060 22204 27580 22260
rect 27636 22204 27646 22260
rect 49970 22204 49980 22260
rect 50036 22204 50988 22260
rect 51044 22204 51054 22260
rect 51426 22204 51436 22260
rect 51492 22204 52668 22260
rect 52724 22204 52734 22260
rect 2930 22092 2940 22148
rect 2996 22092 5964 22148
rect 6020 22092 6030 22148
rect 17714 22092 17724 22148
rect 17780 22092 18620 22148
rect 18676 22092 18686 22148
rect 29474 22092 29484 22148
rect 29540 22092 30380 22148
rect 30436 22092 30828 22148
rect 30884 22092 30894 22148
rect 41570 22092 41580 22148
rect 41636 22092 47180 22148
rect 47236 22092 47246 22148
rect 54200 22036 55000 22064
rect 5282 21980 5292 22036
rect 5348 21980 6076 22036
rect 6132 21980 6142 22036
rect 42466 21980 42476 22036
rect 42532 21980 43708 22036
rect 43764 21980 44044 22036
rect 44100 21980 44110 22036
rect 53218 21980 53228 22036
rect 53284 21980 55000 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 54200 21952 55000 21980
rect 5394 21756 5404 21812
rect 5460 21756 7868 21812
rect 7924 21756 7934 21812
rect 34738 21756 34748 21812
rect 34804 21756 38668 21812
rect 38724 21756 38734 21812
rect 39778 21756 39788 21812
rect 39844 21756 42140 21812
rect 42196 21756 42700 21812
rect 42756 21756 42766 21812
rect 44482 21756 44492 21812
rect 44548 21756 44558 21812
rect 5842 21644 5852 21700
rect 5908 21644 6188 21700
rect 6244 21644 7308 21700
rect 7364 21644 7374 21700
rect 24518 21644 24556 21700
rect 24612 21644 24622 21700
rect 30034 21644 30044 21700
rect 30100 21644 35308 21700
rect 35364 21644 35374 21700
rect 35634 21644 35644 21700
rect 35700 21644 42364 21700
rect 42420 21644 42430 21700
rect 44492 21588 44548 21756
rect 46722 21644 46732 21700
rect 46788 21644 47740 21700
rect 47796 21644 47806 21700
rect 52658 21644 52668 21700
rect 52724 21644 53228 21700
rect 53284 21644 53294 21700
rect 6626 21532 6636 21588
rect 6692 21532 7420 21588
rect 7476 21532 7486 21588
rect 16818 21532 16828 21588
rect 16884 21532 17724 21588
rect 17780 21532 17790 21588
rect 23986 21532 23996 21588
rect 24052 21532 24220 21588
rect 24276 21532 24286 21588
rect 34850 21532 34860 21588
rect 34916 21532 36092 21588
rect 36148 21532 36158 21588
rect 37762 21532 37772 21588
rect 37828 21532 40572 21588
rect 40628 21532 40638 21588
rect 41570 21532 41580 21588
rect 41636 21532 43932 21588
rect 43988 21532 43998 21588
rect 44156 21532 44548 21588
rect 44156 21476 44212 21532
rect 6290 21420 6300 21476
rect 6356 21420 7196 21476
rect 7252 21420 7262 21476
rect 21298 21420 21308 21476
rect 21364 21420 23548 21476
rect 23604 21420 23614 21476
rect 30370 21420 30380 21476
rect 30436 21420 35644 21476
rect 35700 21420 35710 21476
rect 36194 21420 36204 21476
rect 36260 21420 44212 21476
rect 44482 21420 44492 21476
rect 44548 21420 45052 21476
rect 45108 21420 45118 21476
rect 17490 21308 17500 21364
rect 17556 21308 18284 21364
rect 18340 21308 32732 21364
rect 32788 21308 32798 21364
rect 34290 21308 34300 21364
rect 34356 21308 37100 21364
rect 37156 21308 37166 21364
rect 38612 21308 41020 21364
rect 41076 21308 41086 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 7746 21084 7756 21140
rect 7812 21084 11340 21140
rect 11396 21084 11406 21140
rect 38612 21028 38668 21308
rect 41010 21084 41020 21140
rect 41076 21084 43148 21140
rect 43204 21084 43214 21140
rect 33954 20972 33964 21028
rect 34020 20972 38668 21028
rect 42018 20972 42028 21028
rect 42084 20972 42700 21028
rect 42756 20972 42766 21028
rect 11330 20860 11340 20916
rect 11396 20860 25228 20916
rect 25284 20860 29932 20916
rect 29988 20860 29998 20916
rect 32386 20860 32396 20916
rect 32452 20860 32956 20916
rect 33012 20860 37772 20916
rect 37828 20860 37838 20916
rect 41458 20860 41468 20916
rect 41524 20860 43372 20916
rect 43428 20860 43438 20916
rect 37650 20748 37660 20804
rect 37716 20748 39116 20804
rect 39172 20748 39182 20804
rect 40226 20748 40236 20804
rect 40292 20748 42140 20804
rect 42196 20748 42206 20804
rect 45154 20748 45164 20804
rect 45220 20748 45230 20804
rect 45378 20748 45388 20804
rect 45444 20748 45948 20804
rect 46004 20748 46014 20804
rect 45164 20692 45220 20748
rect 9884 20636 16716 20692
rect 16772 20636 16782 20692
rect 29138 20636 29148 20692
rect 29204 20636 30044 20692
rect 30100 20636 30828 20692
rect 30884 20636 30894 20692
rect 35970 20636 35980 20692
rect 36036 20636 37324 20692
rect 37380 20636 37390 20692
rect 41570 20636 41580 20692
rect 41636 20636 44156 20692
rect 44212 20636 44222 20692
rect 45164 20636 46284 20692
rect 46340 20636 46350 20692
rect 3042 20524 3052 20580
rect 3108 20524 5740 20580
rect 5796 20524 5806 20580
rect 9884 20356 9940 20636
rect 11890 20524 11900 20580
rect 11956 20524 16604 20580
rect 16660 20524 16670 20580
rect 18732 20524 31500 20580
rect 31556 20524 31566 20580
rect 32050 20524 32060 20580
rect 32116 20524 33516 20580
rect 33572 20524 41692 20580
rect 41748 20524 41758 20580
rect 49858 20524 49868 20580
rect 49924 20524 51548 20580
rect 51604 20524 51614 20580
rect 18732 20468 18788 20524
rect 16034 20412 16044 20468
rect 16100 20412 18788 20468
rect 44230 20412 44268 20468
rect 44324 20412 44334 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 9874 20300 9884 20356
rect 9940 20300 9950 20356
rect 24098 20300 24108 20356
rect 24164 20300 26796 20356
rect 26852 20300 26862 20356
rect 44146 20300 44156 20356
rect 44212 20300 44772 20356
rect 44930 20300 44940 20356
rect 44996 20300 45500 20356
rect 45556 20300 45566 20356
rect 1698 20188 1708 20244
rect 1764 20188 4844 20244
rect 4900 20188 9660 20244
rect 9716 20188 9726 20244
rect 10546 20188 10556 20244
rect 10612 20188 11340 20244
rect 11396 20188 11406 20244
rect 39890 20188 39900 20244
rect 39956 20188 40236 20244
rect 40292 20188 40302 20244
rect 42466 20188 42476 20244
rect 42532 20188 43932 20244
rect 43988 20188 44492 20244
rect 44548 20188 44558 20244
rect 44716 20132 44772 20300
rect 45378 20188 45388 20244
rect 45444 20188 46732 20244
rect 46788 20188 46798 20244
rect 50306 20188 50316 20244
rect 50372 20188 50382 20244
rect 50316 20132 50372 20188
rect 2818 20076 2828 20132
rect 2884 20076 3500 20132
rect 3556 20076 3566 20132
rect 11778 20076 11788 20132
rect 11844 20076 13020 20132
rect 13076 20076 14700 20132
rect 14756 20076 14766 20132
rect 15026 20076 15036 20132
rect 15092 20076 15708 20132
rect 15764 20076 31836 20132
rect 31892 20076 31902 20132
rect 33170 20076 33180 20132
rect 33236 20076 34300 20132
rect 34356 20076 34366 20132
rect 39218 20076 39228 20132
rect 39284 20076 41132 20132
rect 41188 20076 41580 20132
rect 41636 20076 41646 20132
rect 41794 20076 41804 20132
rect 41860 20076 42812 20132
rect 42868 20076 45052 20132
rect 45108 20076 45118 20132
rect 46834 20076 46844 20132
rect 46900 20076 47516 20132
rect 47572 20076 47582 20132
rect 49756 20076 50372 20132
rect 3332 19460 3388 20076
rect 49756 20020 49812 20076
rect 4946 19964 4956 20020
rect 5012 19964 5180 20020
rect 5236 19964 5628 20020
rect 5684 19964 15484 20020
rect 15540 19964 15550 20020
rect 24770 19964 24780 20020
rect 24836 19964 26124 20020
rect 26180 19964 26572 20020
rect 26628 19964 26638 20020
rect 30258 19964 30268 20020
rect 30324 19964 30828 20020
rect 30884 19964 30894 20020
rect 32162 19964 32172 20020
rect 32228 19964 33068 20020
rect 33124 19964 33134 20020
rect 34738 19964 34748 20020
rect 34804 19964 38668 20020
rect 39442 19964 39452 20020
rect 39508 19964 39788 20020
rect 39844 19964 39854 20020
rect 41458 19964 41468 20020
rect 41524 19964 42140 20020
rect 42196 19964 42206 20020
rect 44482 19964 44492 20020
rect 44548 19964 45612 20020
rect 45668 19964 47292 20020
rect 47348 19964 47358 20020
rect 48066 19964 48076 20020
rect 48132 19964 49756 20020
rect 49812 19964 49822 20020
rect 38612 19908 38668 19964
rect 8082 19852 8092 19908
rect 8148 19852 8652 19908
rect 8708 19852 9324 19908
rect 9380 19852 16044 19908
rect 16100 19852 16110 19908
rect 16258 19852 16268 19908
rect 16324 19852 17500 19908
rect 17556 19852 17566 19908
rect 21410 19852 21420 19908
rect 21476 19852 23884 19908
rect 23940 19852 23950 19908
rect 29474 19852 29484 19908
rect 29540 19852 37100 19908
rect 37156 19852 37166 19908
rect 38612 19852 43708 19908
rect 43764 19852 44604 19908
rect 44660 19852 46060 19908
rect 46116 19852 46126 19908
rect 51314 19852 51324 19908
rect 51380 19852 51772 19908
rect 51828 19852 53228 19908
rect 53284 19852 53294 19908
rect 7074 19740 7084 19796
rect 7140 19740 8204 19796
rect 8260 19740 10220 19796
rect 10276 19740 10286 19796
rect 20514 19740 20524 19796
rect 20580 19740 30492 19796
rect 30548 19740 31388 19796
rect 31444 19740 31454 19796
rect 47842 19740 47852 19796
rect 47908 19740 48748 19796
rect 48804 19740 48814 19796
rect 20290 19628 20300 19684
rect 20356 19628 32844 19684
rect 32900 19628 32910 19684
rect 44146 19628 44156 19684
rect 44212 19628 44940 19684
rect 44996 19628 45006 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 3332 19404 20412 19460
rect 20468 19404 20478 19460
rect 23090 19404 23100 19460
rect 23156 19404 23548 19460
rect 26562 19404 26572 19460
rect 26628 19404 37772 19460
rect 37828 19404 37838 19460
rect 44230 19404 44268 19460
rect 44324 19404 44334 19460
rect 9538 19292 9548 19348
rect 9604 19292 17052 19348
rect 17108 19292 18172 19348
rect 18228 19292 18238 19348
rect 7522 19068 7532 19124
rect 7588 19068 11452 19124
rect 11508 19068 11518 19124
rect 23492 19012 23548 19404
rect 54200 19348 55000 19376
rect 24098 19292 24108 19348
rect 24164 19292 24444 19348
rect 24500 19292 24510 19348
rect 32722 19292 32732 19348
rect 32788 19292 45836 19348
rect 45892 19292 45902 19348
rect 49298 19292 49308 19348
rect 49364 19292 50316 19348
rect 50372 19292 50382 19348
rect 52210 19292 52220 19348
rect 52276 19292 53228 19348
rect 53284 19292 55000 19348
rect 54200 19264 55000 19292
rect 23958 19180 23996 19236
rect 24052 19180 24062 19236
rect 24546 19180 24556 19236
rect 24612 19180 25340 19236
rect 25396 19180 25406 19236
rect 29362 19180 29372 19236
rect 29428 19180 30268 19236
rect 30324 19180 30334 19236
rect 32498 19180 32508 19236
rect 32564 19180 33628 19236
rect 33684 19180 34524 19236
rect 34580 19180 34590 19236
rect 41234 19180 41244 19236
rect 41300 19180 41692 19236
rect 41748 19180 41758 19236
rect 43810 19180 43820 19236
rect 43876 19180 45444 19236
rect 28466 19068 28476 19124
rect 28532 19068 29316 19124
rect 33394 19068 33404 19124
rect 33460 19068 39564 19124
rect 39620 19068 41356 19124
rect 41412 19068 41916 19124
rect 41972 19068 43484 19124
rect 43540 19068 43550 19124
rect 29260 19012 29316 19068
rect 45388 19012 45444 19180
rect 47730 19068 47740 19124
rect 47796 19068 49084 19124
rect 49140 19068 49150 19124
rect 20178 18956 20188 19012
rect 20244 18956 23324 19012
rect 23380 18956 23390 19012
rect 23492 18956 24332 19012
rect 24388 18956 24398 19012
rect 27570 18956 27580 19012
rect 27636 18956 29036 19012
rect 29092 18956 29102 19012
rect 29250 18956 29260 19012
rect 29316 18956 29820 19012
rect 29876 18956 36428 19012
rect 36484 18956 38780 19012
rect 38836 18956 38846 19012
rect 42354 18956 42364 19012
rect 42420 18956 44268 19012
rect 44324 18956 44334 19012
rect 45378 18956 45388 19012
rect 45444 18956 46396 19012
rect 46452 18956 46462 19012
rect 31266 18844 31276 18900
rect 31332 18844 31836 18900
rect 31892 18844 33740 18900
rect 33796 18844 34300 18900
rect 34356 18844 38668 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 31490 18620 31500 18676
rect 31556 18620 34076 18676
rect 34132 18620 34142 18676
rect 38612 18564 38668 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 6850 18508 6860 18564
rect 6916 18508 7532 18564
rect 7588 18508 7598 18564
rect 14466 18508 14476 18564
rect 14532 18508 15372 18564
rect 15428 18508 15438 18564
rect 25106 18508 25116 18564
rect 25172 18508 26572 18564
rect 26628 18508 27132 18564
rect 27188 18508 27198 18564
rect 31938 18508 31948 18564
rect 32004 18508 32508 18564
rect 32564 18508 32574 18564
rect 38612 18508 42868 18564
rect 6626 18396 6636 18452
rect 6692 18396 7980 18452
rect 8036 18396 8046 18452
rect 8306 18396 8316 18452
rect 8372 18396 8988 18452
rect 9044 18396 9772 18452
rect 9828 18396 9838 18452
rect 12562 18396 12572 18452
rect 12628 18396 13580 18452
rect 13636 18396 16268 18452
rect 16324 18396 16334 18452
rect 26226 18396 26236 18452
rect 26292 18396 27020 18452
rect 27076 18396 27086 18452
rect 31490 18396 31500 18452
rect 31556 18396 32172 18452
rect 32228 18396 32238 18452
rect 40338 18396 40348 18452
rect 40404 18396 40908 18452
rect 40964 18396 42588 18452
rect 42644 18396 42654 18452
rect 7196 18228 7252 18396
rect 42812 18340 42868 18508
rect 43138 18396 43148 18452
rect 43204 18396 50988 18452
rect 51044 18396 51054 18452
rect 51874 18396 51884 18452
rect 51940 18396 52444 18452
rect 52500 18396 52510 18452
rect 15922 18284 15932 18340
rect 15988 18284 24892 18340
rect 24948 18284 24958 18340
rect 29922 18284 29932 18340
rect 29988 18284 31612 18340
rect 31668 18284 31678 18340
rect 42812 18284 44492 18340
rect 44548 18284 44558 18340
rect 46274 18284 46284 18340
rect 46340 18284 48636 18340
rect 48692 18284 49644 18340
rect 49700 18284 49710 18340
rect 7186 18172 7196 18228
rect 7252 18172 7262 18228
rect 43810 18172 43820 18228
rect 43876 18172 48748 18228
rect 48804 18172 48814 18228
rect 51212 18172 52220 18228
rect 52276 18172 52286 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 51212 18004 51268 18172
rect 23426 17948 23436 18004
rect 23492 17948 31836 18004
rect 31892 17948 31902 18004
rect 51202 17948 51212 18004
rect 51268 17948 51278 18004
rect 51762 17948 51772 18004
rect 51828 17948 52108 18004
rect 52164 17948 52174 18004
rect 9650 17836 9660 17892
rect 9716 17836 9726 17892
rect 31714 17836 31724 17892
rect 31780 17836 32620 17892
rect 32676 17836 38892 17892
rect 38948 17836 38958 17892
rect 9660 17780 9716 17836
rect 9090 17724 9100 17780
rect 9156 17724 10108 17780
rect 10164 17724 10668 17780
rect 10724 17724 14364 17780
rect 14420 17724 14430 17780
rect 33170 17724 33180 17780
rect 33236 17724 35420 17780
rect 35476 17724 36540 17780
rect 36596 17724 40684 17780
rect 40740 17724 40750 17780
rect 45154 17724 45164 17780
rect 45220 17724 50428 17780
rect 6178 17612 6188 17668
rect 6244 17612 7420 17668
rect 7476 17612 9660 17668
rect 9716 17612 9726 17668
rect 32386 17612 32396 17668
rect 32452 17612 33068 17668
rect 33124 17612 33134 17668
rect 38994 17612 39004 17668
rect 39060 17612 40572 17668
rect 40628 17612 40638 17668
rect 45938 17612 45948 17668
rect 46004 17612 49196 17668
rect 49252 17612 49262 17668
rect 50372 17556 50428 17724
rect 50978 17612 50988 17668
rect 51044 17612 51212 17668
rect 51268 17612 53004 17668
rect 53060 17612 53070 17668
rect 24322 17500 24332 17556
rect 24388 17500 24668 17556
rect 24724 17500 25788 17556
rect 25844 17500 25854 17556
rect 38210 17500 38220 17556
rect 38276 17500 39228 17556
rect 39284 17500 39294 17556
rect 44146 17500 44156 17556
rect 44212 17500 45500 17556
rect 45556 17500 45566 17556
rect 50372 17500 50652 17556
rect 50708 17500 52780 17556
rect 52836 17500 52846 17556
rect 6738 17388 6748 17444
rect 6804 17388 8316 17444
rect 8372 17388 8382 17444
rect 16370 17388 16380 17444
rect 16436 17388 17052 17444
rect 17108 17388 22764 17444
rect 22820 17388 22830 17444
rect 25666 17388 25676 17444
rect 25732 17388 28252 17444
rect 28308 17388 28318 17444
rect 34178 17388 34188 17444
rect 34244 17388 36428 17444
rect 36484 17388 37548 17444
rect 37604 17388 37614 17444
rect 38546 17388 38556 17444
rect 38612 17388 39564 17444
rect 39620 17388 43148 17444
rect 43204 17388 47852 17444
rect 47908 17388 47918 17444
rect 49186 17388 49196 17444
rect 49252 17388 50540 17444
rect 50596 17388 51100 17444
rect 51156 17388 51166 17444
rect 51874 17388 51884 17444
rect 51940 17388 52556 17444
rect 52612 17388 52622 17444
rect 33170 17276 33180 17332
rect 33236 17276 44604 17332
rect 44660 17276 44670 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 15474 17164 15484 17220
rect 15540 17164 17612 17220
rect 17668 17164 17678 17220
rect 32722 17164 32732 17220
rect 32788 17164 36652 17220
rect 36708 17164 38668 17220
rect 38724 17164 38734 17220
rect 40226 17164 40236 17220
rect 40292 17164 41244 17220
rect 41300 17164 41310 17220
rect 42578 17164 42588 17220
rect 42644 17164 43932 17220
rect 43988 17164 44940 17220
rect 44996 17164 45006 17220
rect 46274 17164 46284 17220
rect 46340 17164 47404 17220
rect 47460 17164 47470 17220
rect 2482 17052 2492 17108
rect 2548 17052 6412 17108
rect 6468 17052 6478 17108
rect 14802 17052 14812 17108
rect 14868 17052 15820 17108
rect 15876 17052 15886 17108
rect 16482 17052 16492 17108
rect 16548 17052 17948 17108
rect 18004 17052 18014 17108
rect 23762 17052 23772 17108
rect 23828 17052 24220 17108
rect 24276 17052 24556 17108
rect 24612 17052 24622 17108
rect 30258 17052 30268 17108
rect 30324 17052 37996 17108
rect 38052 17052 38556 17108
rect 38612 17052 38622 17108
rect 42914 17052 42924 17108
rect 42980 17052 51324 17108
rect 51380 17052 51772 17108
rect 51828 17052 51838 17108
rect 13906 16940 13916 16996
rect 13972 16940 15652 16996
rect 38658 16940 38668 16996
rect 38724 16940 40236 16996
rect 40292 16940 40302 16996
rect 45042 16940 45052 16996
rect 45108 16940 49308 16996
rect 49364 16940 52892 16996
rect 52948 16940 52958 16996
rect 15596 16884 15652 16940
rect 6850 16828 6860 16884
rect 6916 16828 7532 16884
rect 7588 16828 7598 16884
rect 11106 16828 11116 16884
rect 11172 16828 11900 16884
rect 11956 16828 13132 16884
rect 13188 16828 13198 16884
rect 13458 16828 13468 16884
rect 13524 16828 14588 16884
rect 14644 16828 14654 16884
rect 15596 16828 17276 16884
rect 17332 16828 17342 16884
rect 17490 16828 17500 16884
rect 17556 16828 20076 16884
rect 20132 16828 20142 16884
rect 34178 16828 34188 16884
rect 34244 16828 38108 16884
rect 38164 16828 39004 16884
rect 39060 16828 39070 16884
rect 39442 16828 39452 16884
rect 39508 16828 41020 16884
rect 41076 16828 41086 16884
rect 45490 16828 45500 16884
rect 45556 16828 46844 16884
rect 46900 16828 46910 16884
rect 52658 16828 52668 16884
rect 52724 16828 53228 16884
rect 53284 16828 53294 16884
rect 16146 16716 16156 16772
rect 16212 16716 17836 16772
rect 17892 16716 17902 16772
rect 19058 16716 19068 16772
rect 19124 16716 21084 16772
rect 21140 16716 21150 16772
rect 21634 16716 21644 16772
rect 21700 16716 23324 16772
rect 23380 16716 23390 16772
rect 24098 16716 24108 16772
rect 24164 16716 24892 16772
rect 24948 16716 25228 16772
rect 25284 16716 25294 16772
rect 35970 16716 35980 16772
rect 36036 16716 36316 16772
rect 36372 16716 39340 16772
rect 39396 16716 39406 16772
rect 42578 16716 42588 16772
rect 42644 16716 44156 16772
rect 44212 16716 44222 16772
rect 53228 16660 53284 16828
rect 54200 16660 55000 16688
rect 14914 16604 14924 16660
rect 14980 16604 16492 16660
rect 16548 16604 16558 16660
rect 44258 16604 44268 16660
rect 44324 16604 51548 16660
rect 51604 16604 51614 16660
rect 53228 16604 55000 16660
rect 54200 16576 55000 16604
rect 4946 16492 4956 16548
rect 5012 16492 5628 16548
rect 5684 16492 6300 16548
rect 6356 16492 6636 16548
rect 6692 16492 6702 16548
rect 38322 16492 38332 16548
rect 38388 16492 39564 16548
rect 39620 16492 39630 16548
rect 46610 16492 46620 16548
rect 46676 16492 49196 16548
rect 49252 16492 49262 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 50866 16380 50876 16436
rect 50932 16380 50942 16436
rect 12898 16268 12908 16324
rect 12964 16268 13580 16324
rect 13636 16268 13646 16324
rect 16594 16268 16604 16324
rect 16660 16268 17388 16324
rect 17444 16268 17454 16324
rect 40338 16268 40348 16324
rect 40404 16268 43820 16324
rect 43876 16268 44716 16324
rect 44772 16268 44782 16324
rect 4610 16156 4620 16212
rect 4676 16156 5404 16212
rect 5460 16156 6188 16212
rect 6244 16156 6254 16212
rect 40226 16156 40236 16212
rect 40292 16156 44268 16212
rect 44324 16156 44334 16212
rect 5282 16044 5292 16100
rect 5348 16044 9660 16100
rect 9716 16044 13580 16100
rect 13636 16044 16716 16100
rect 16772 16044 16782 16100
rect 23090 16044 23100 16100
rect 23156 16044 25116 16100
rect 25172 16044 25182 16100
rect 38994 16044 39004 16100
rect 39060 16044 42364 16100
rect 42420 16044 42430 16100
rect 5058 15932 5068 15988
rect 5124 15932 5964 15988
rect 6020 15932 6030 15988
rect 15810 15932 15820 15988
rect 15876 15932 16044 15988
rect 16100 15932 17276 15988
rect 17332 15932 17342 15988
rect 24434 15932 24444 15988
rect 24500 15932 28812 15988
rect 28868 15932 28878 15988
rect 39218 15932 39228 15988
rect 39284 15932 39788 15988
rect 39844 15932 39854 15988
rect 40012 15876 40068 16044
rect 50876 15988 50932 16380
rect 49186 15932 49196 15988
rect 49252 15932 49756 15988
rect 49812 15932 49822 15988
rect 49970 15932 49980 15988
rect 50036 15932 50428 15988
rect 50484 15932 50494 15988
rect 50876 15932 52668 15988
rect 52724 15932 52734 15988
rect 10210 15820 10220 15876
rect 10276 15820 13580 15876
rect 13636 15820 14252 15876
rect 14308 15820 14318 15876
rect 34290 15820 34300 15876
rect 34356 15820 36204 15876
rect 36260 15820 37660 15876
rect 37716 15820 37726 15876
rect 39554 15820 39564 15876
rect 39620 15820 40068 15876
rect 50642 15820 50652 15876
rect 50708 15820 51324 15876
rect 51380 15820 51390 15876
rect 51762 15820 51772 15876
rect 51828 15820 52780 15876
rect 52836 15820 52846 15876
rect 25330 15708 25340 15764
rect 25396 15708 29260 15764
rect 29316 15708 29326 15764
rect 38546 15708 38556 15764
rect 38612 15708 40348 15764
rect 40404 15708 40414 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 6514 15484 6524 15540
rect 6580 15484 10332 15540
rect 10388 15484 10398 15540
rect 18162 15484 18172 15540
rect 18228 15484 19516 15540
rect 19572 15484 19582 15540
rect 35298 15484 35308 15540
rect 35364 15484 36428 15540
rect 36484 15484 36494 15540
rect 45490 15484 45500 15540
rect 45556 15484 46172 15540
rect 46228 15484 46238 15540
rect 49074 15484 49084 15540
rect 49140 15484 49644 15540
rect 49700 15484 49710 15540
rect 49868 15484 50316 15540
rect 50372 15484 52332 15540
rect 52388 15484 52398 15540
rect 45500 15428 45556 15484
rect 6066 15372 6076 15428
rect 6132 15372 8652 15428
rect 8708 15372 8718 15428
rect 10546 15372 10556 15428
rect 10612 15372 12908 15428
rect 12964 15372 12974 15428
rect 38612 15372 38780 15428
rect 38836 15372 38846 15428
rect 42690 15372 42700 15428
rect 42756 15372 45556 15428
rect 11218 15260 11228 15316
rect 11284 15260 14588 15316
rect 14644 15260 14654 15316
rect 18834 15260 18844 15316
rect 18900 15260 20972 15316
rect 21028 15260 22092 15316
rect 22148 15260 24108 15316
rect 24164 15260 28476 15316
rect 28532 15260 29596 15316
rect 29652 15260 29662 15316
rect 32050 15260 32060 15316
rect 32116 15260 33796 15316
rect 35634 15260 35644 15316
rect 35700 15260 37324 15316
rect 37380 15260 37390 15316
rect 33740 15204 33796 15260
rect 38612 15204 38668 15372
rect 49868 15316 49924 15484
rect 50082 15372 50092 15428
rect 50148 15372 53116 15428
rect 53172 15372 53182 15428
rect 45266 15260 45276 15316
rect 45332 15260 45836 15316
rect 45892 15260 46284 15316
rect 46340 15260 46350 15316
rect 46498 15260 46508 15316
rect 46564 15260 49084 15316
rect 49140 15260 49924 15316
rect 50372 15260 51100 15316
rect 51156 15260 51166 15316
rect 50372 15204 50428 15260
rect 32498 15148 32508 15204
rect 32564 15148 33404 15204
rect 33460 15148 33470 15204
rect 33730 15148 33740 15204
rect 33796 15148 38668 15204
rect 42466 15148 42476 15204
rect 42532 15148 43484 15204
rect 43540 15148 43550 15204
rect 48626 15148 48636 15204
rect 48692 15148 50428 15204
rect 51314 15148 51324 15204
rect 51380 15148 52108 15204
rect 52164 15148 52174 15204
rect 6402 15036 6412 15092
rect 6468 15036 6860 15092
rect 6916 15036 8092 15092
rect 8148 15036 8158 15092
rect 20290 15036 20300 15092
rect 20356 15036 47628 15092
rect 47684 15036 52668 15092
rect 52724 15036 52734 15092
rect 26786 14924 26796 14980
rect 26852 14924 27580 14980
rect 27636 14924 31164 14980
rect 31220 14924 31230 14980
rect 44146 14924 44156 14980
rect 44212 14924 44716 14980
rect 44772 14924 44782 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 29474 14812 29484 14868
rect 29540 14812 31052 14868
rect 31108 14812 31118 14868
rect 6626 14700 6636 14756
rect 6692 14700 8316 14756
rect 8372 14700 8382 14756
rect 45378 14700 45388 14756
rect 45444 14700 45948 14756
rect 46004 14700 46014 14756
rect 9202 14588 9212 14644
rect 9268 14588 9660 14644
rect 9716 14588 10108 14644
rect 10164 14588 10174 14644
rect 30146 14588 30156 14644
rect 30212 14588 40908 14644
rect 40964 14588 40974 14644
rect 45826 14588 45836 14644
rect 45892 14588 50204 14644
rect 50260 14588 50270 14644
rect 13010 14476 13020 14532
rect 13076 14476 15148 14532
rect 15204 14476 15708 14532
rect 15764 14476 15774 14532
rect 17378 14476 17388 14532
rect 17444 14476 19068 14532
rect 19124 14476 19134 14532
rect 24322 14476 24332 14532
rect 24388 14476 24668 14532
rect 24724 14476 26012 14532
rect 26068 14476 26078 14532
rect 38210 14476 38220 14532
rect 38276 14476 46284 14532
rect 46340 14476 46350 14532
rect 15362 14364 15372 14420
rect 15428 14364 16380 14420
rect 16436 14364 17164 14420
rect 17220 14364 17230 14420
rect 17714 14364 17724 14420
rect 17780 14364 18396 14420
rect 18452 14364 18462 14420
rect 38434 14364 38444 14420
rect 38500 14364 39676 14420
rect 39732 14364 39742 14420
rect 40114 14364 40124 14420
rect 40180 14364 41916 14420
rect 41972 14364 41982 14420
rect 43922 14364 43932 14420
rect 43988 14364 52668 14420
rect 52724 14364 52734 14420
rect 8194 14252 8204 14308
rect 8260 14252 8876 14308
rect 8932 14252 8942 14308
rect 16034 14252 16044 14308
rect 16100 14252 18284 14308
rect 18340 14252 18350 14308
rect 24210 14252 24220 14308
rect 24276 14252 25340 14308
rect 25396 14252 25406 14308
rect 26114 14252 26124 14308
rect 26180 14252 29484 14308
rect 29540 14252 29550 14308
rect 30706 14252 30716 14308
rect 30772 14252 31500 14308
rect 31556 14252 31566 14308
rect 47394 14252 47404 14308
rect 47460 14252 48524 14308
rect 48580 14252 52892 14308
rect 52948 14252 52958 14308
rect 8754 14140 8764 14196
rect 8820 14140 9436 14196
rect 9492 14140 9502 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 10098 14028 10108 14084
rect 10164 14028 10780 14084
rect 10836 14028 11564 14084
rect 11620 14028 13132 14084
rect 13188 14028 13198 14084
rect 54200 13972 55000 14000
rect 6626 13916 6636 13972
rect 6692 13916 7420 13972
rect 7476 13916 7486 13972
rect 11890 13916 11900 13972
rect 11956 13916 46844 13972
rect 46900 13916 46910 13972
rect 53330 13916 53340 13972
rect 53396 13916 55000 13972
rect 54200 13888 55000 13916
rect 7522 13804 7532 13860
rect 7588 13804 9212 13860
rect 9268 13804 12348 13860
rect 12404 13804 14364 13860
rect 14420 13804 14430 13860
rect 35970 13804 35980 13860
rect 36036 13804 39004 13860
rect 39060 13804 40124 13860
rect 40180 13804 41356 13860
rect 41412 13804 41422 13860
rect 4946 13692 4956 13748
rect 5012 13692 5628 13748
rect 5684 13692 5694 13748
rect 8082 13692 8092 13748
rect 8148 13692 8652 13748
rect 8708 13692 8718 13748
rect 24658 13692 24668 13748
rect 24724 13692 26572 13748
rect 26628 13692 26638 13748
rect 36642 13692 36652 13748
rect 36708 13692 39676 13748
rect 39732 13692 39742 13748
rect 46358 13692 46396 13748
rect 46452 13692 46462 13748
rect 21746 13580 21756 13636
rect 21812 13580 24220 13636
rect 24276 13580 24286 13636
rect 24434 13580 24444 13636
rect 24500 13580 25340 13636
rect 25396 13580 25788 13636
rect 25844 13580 25854 13636
rect 26114 13580 26124 13636
rect 26180 13580 27356 13636
rect 27412 13580 27422 13636
rect 39106 13580 39116 13636
rect 39172 13580 40908 13636
rect 40964 13580 41804 13636
rect 41860 13580 41870 13636
rect 42578 13580 42588 13636
rect 42644 13580 43932 13636
rect 43988 13580 43998 13636
rect 17938 13468 17948 13524
rect 18004 13468 18508 13524
rect 18564 13468 20860 13524
rect 20916 13468 20926 13524
rect 44594 13468 44604 13524
rect 44660 13468 45948 13524
rect 46004 13468 46732 13524
rect 46788 13468 46798 13524
rect 48178 13468 48188 13524
rect 48244 13468 49196 13524
rect 49252 13468 50372 13524
rect 51090 13468 51100 13524
rect 51156 13468 52220 13524
rect 52276 13468 52286 13524
rect 50316 13412 50372 13468
rect 6850 13356 6860 13412
rect 6916 13356 7644 13412
rect 7700 13356 7710 13412
rect 14130 13356 14140 13412
rect 14196 13356 14588 13412
rect 14644 13356 23436 13412
rect 23492 13356 23502 13412
rect 40198 13356 40236 13412
rect 40292 13356 40302 13412
rect 41794 13356 41804 13412
rect 41860 13356 45388 13412
rect 45444 13356 45454 13412
rect 50306 13356 50316 13412
rect 50372 13356 51436 13412
rect 51492 13356 51502 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 26674 13244 26684 13300
rect 26740 13244 27020 13300
rect 27076 13244 27086 13300
rect 29362 13244 29372 13300
rect 29428 13244 35028 13300
rect 34972 13188 35028 13244
rect 13906 13132 13916 13188
rect 13972 13132 15932 13188
rect 15988 13132 17612 13188
rect 17668 13132 17678 13188
rect 19058 13132 19068 13188
rect 19124 13132 30156 13188
rect 30212 13132 30222 13188
rect 30380 13132 33180 13188
rect 33236 13132 33246 13188
rect 34972 13132 37548 13188
rect 37604 13132 37614 13188
rect 19068 13076 19124 13132
rect 30380 13076 30436 13132
rect 17378 13020 17388 13076
rect 17444 13020 19124 13076
rect 19964 13020 30436 13076
rect 31826 13020 31836 13076
rect 31892 13020 31902 13076
rect 35634 13020 35644 13076
rect 35700 13020 35710 13076
rect 42466 13020 42476 13076
rect 42532 13020 43036 13076
rect 43092 13020 45836 13076
rect 45892 13020 45902 13076
rect 2594 12908 2604 12964
rect 2660 12908 8204 12964
rect 8260 12908 8270 12964
rect 17826 12908 17836 12964
rect 17892 12908 18396 12964
rect 18452 12908 18462 12964
rect 19964 12852 20020 13020
rect 31836 12852 31892 13020
rect 35644 12964 35700 13020
rect 33618 12908 33628 12964
rect 33684 12908 34748 12964
rect 34804 12908 37436 12964
rect 37492 12908 37502 12964
rect 38322 12908 38332 12964
rect 38388 12908 39116 12964
rect 39172 12908 39182 12964
rect 41010 12908 41020 12964
rect 41076 12908 42252 12964
rect 42308 12908 42318 12964
rect 7868 12796 8428 12852
rect 8484 12796 9100 12852
rect 9156 12796 9166 12852
rect 16146 12796 16156 12852
rect 16212 12796 16828 12852
rect 16884 12796 20020 12852
rect 26114 12796 26124 12852
rect 26180 12796 27132 12852
rect 27188 12796 27198 12852
rect 31836 12796 36092 12852
rect 36148 12796 36158 12852
rect 39554 12796 39564 12852
rect 39620 12796 40460 12852
rect 40516 12796 40526 12852
rect 7868 12516 7924 12796
rect 11218 12684 11228 12740
rect 11284 12684 13468 12740
rect 13524 12684 13534 12740
rect 15138 12684 15148 12740
rect 15204 12684 16044 12740
rect 16100 12684 16110 12740
rect 22866 12684 22876 12740
rect 22932 12684 26572 12740
rect 26628 12684 26638 12740
rect 35634 12684 35644 12740
rect 35700 12684 36204 12740
rect 36260 12684 36270 12740
rect 36418 12684 36428 12740
rect 36484 12684 38108 12740
rect 38164 12684 38174 12740
rect 15250 12572 15260 12628
rect 15316 12572 15326 12628
rect 34850 12572 34860 12628
rect 34916 12572 34926 12628
rect 15260 12516 15316 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 5282 12460 5292 12516
rect 5348 12460 5740 12516
rect 5796 12460 7868 12516
rect 7924 12460 7934 12516
rect 15148 12460 15316 12516
rect 6850 12348 6860 12404
rect 6916 12348 8428 12404
rect 8484 12348 8494 12404
rect 7410 12124 7420 12180
rect 7476 12124 7486 12180
rect 7420 12068 7476 12124
rect 15148 12068 15204 12460
rect 34860 12404 34916 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 27122 12348 27132 12404
rect 27188 12348 28252 12404
rect 28308 12348 30268 12404
rect 30324 12348 30334 12404
rect 34748 12348 35980 12404
rect 36036 12348 36046 12404
rect 16370 12236 16380 12292
rect 16436 12236 18060 12292
rect 18116 12236 18126 12292
rect 23538 12236 23548 12292
rect 23604 12236 24444 12292
rect 24500 12236 24510 12292
rect 34748 12180 34804 12348
rect 38612 12292 38668 12404
rect 38724 12348 38734 12404
rect 36306 12236 36316 12292
rect 36372 12236 37996 12292
rect 38052 12236 38668 12292
rect 15810 12124 15820 12180
rect 15876 12124 18620 12180
rect 18676 12124 18686 12180
rect 23762 12124 23772 12180
rect 23828 12124 24332 12180
rect 24388 12124 24398 12180
rect 24658 12124 24668 12180
rect 24724 12124 25900 12180
rect 25956 12124 25966 12180
rect 33842 12124 33852 12180
rect 33908 12124 34748 12180
rect 34804 12124 34814 12180
rect 38098 12124 38108 12180
rect 38164 12124 38780 12180
rect 38836 12124 38846 12180
rect 45714 12124 45724 12180
rect 45780 12124 49084 12180
rect 49140 12124 49532 12180
rect 49588 12124 49598 12180
rect 2482 12012 2492 12068
rect 2548 12012 6524 12068
rect 6580 12012 6590 12068
rect 7420 12012 8988 12068
rect 9044 12012 9054 12068
rect 15138 12012 15148 12068
rect 15204 12012 15214 12068
rect 23958 12012 23996 12068
rect 24052 12012 24062 12068
rect 26898 12012 26908 12068
rect 26964 12012 30716 12068
rect 30772 12012 30782 12068
rect 35186 12012 35196 12068
rect 35252 12012 39004 12068
rect 39060 12012 40124 12068
rect 40180 12012 41020 12068
rect 41076 12012 41086 12068
rect 41580 12012 42700 12068
rect 42756 12012 42766 12068
rect 51986 12012 51996 12068
rect 52052 12012 53228 12068
rect 53284 12012 53294 12068
rect 41580 11956 41636 12012
rect 6402 11900 6412 11956
rect 6468 11900 7644 11956
rect 7700 11900 7710 11956
rect 23762 11900 23772 11956
rect 23828 11900 25228 11956
rect 25284 11900 25294 11956
rect 37874 11900 37884 11956
rect 37940 11900 41636 11956
rect 21868 11788 25788 11844
rect 25844 11788 25854 11844
rect 26114 11788 26124 11844
rect 26180 11788 26684 11844
rect 26740 11788 26750 11844
rect 38994 11788 39004 11844
rect 39060 11788 39900 11844
rect 39956 11788 40684 11844
rect 40740 11788 40750 11844
rect 40908 11788 42924 11844
rect 42980 11788 42990 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 21868 11732 21924 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 40908 11732 40964 11788
rect 17714 11676 17724 11732
rect 17780 11676 21924 11732
rect 37314 11676 37324 11732
rect 37380 11676 40964 11732
rect 4610 11564 4620 11620
rect 4676 11564 6188 11620
rect 6244 11564 6254 11620
rect 9314 11564 9324 11620
rect 9380 11564 11116 11620
rect 11172 11564 11182 11620
rect 14018 11564 14028 11620
rect 14084 11564 15036 11620
rect 15092 11564 20300 11620
rect 20356 11564 20366 11620
rect 29474 11564 29484 11620
rect 29540 11564 36428 11620
rect 36484 11564 36494 11620
rect 5394 11452 5404 11508
rect 5460 11452 6412 11508
rect 6468 11452 6478 11508
rect 12786 11340 12796 11396
rect 12852 11340 13468 11396
rect 13524 11340 13534 11396
rect 27010 11340 27020 11396
rect 27076 11340 29260 11396
rect 29316 11340 29326 11396
rect 31602 11340 31612 11396
rect 31668 11340 31948 11396
rect 32004 11340 32620 11396
rect 32676 11340 34300 11396
rect 34356 11340 34366 11396
rect 41570 11340 41580 11396
rect 41636 11340 42028 11396
rect 42084 11340 42094 11396
rect 54200 11284 55000 11312
rect 6290 11228 6300 11284
rect 6356 11228 10332 11284
rect 10388 11228 10668 11284
rect 10724 11228 10734 11284
rect 26338 11228 26348 11284
rect 26404 11228 26796 11284
rect 26852 11228 26862 11284
rect 32834 11228 32844 11284
rect 32900 11228 35084 11284
rect 35140 11228 35150 11284
rect 45938 11228 45948 11284
rect 46004 11228 46844 11284
rect 46900 11228 46910 11284
rect 52210 11228 52220 11284
rect 52276 11228 53228 11284
rect 53284 11228 55000 11284
rect 54200 11200 55000 11228
rect 1810 11116 1820 11172
rect 1876 11116 5068 11172
rect 5124 11116 15820 11172
rect 15876 11116 19628 11172
rect 19684 11116 19694 11172
rect 32386 11116 32396 11172
rect 32452 11116 33404 11172
rect 33460 11116 33470 11172
rect 41010 11116 41020 11172
rect 41076 11116 42140 11172
rect 42196 11116 42206 11172
rect 44930 11116 44940 11172
rect 44996 11116 45612 11172
rect 45668 11116 45678 11172
rect 46274 11116 46284 11172
rect 46340 11116 49196 11172
rect 49252 11116 49532 11172
rect 49588 11116 49598 11172
rect 50372 11116 50652 11172
rect 50708 11116 50718 11172
rect 41682 11004 41692 11060
rect 41748 11004 41916 11060
rect 41972 11004 43372 11060
rect 43428 11004 44828 11060
rect 44884 11004 45164 11060
rect 45220 11004 45230 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 30370 10892 30380 10948
rect 30436 10892 35644 10948
rect 35700 10892 41020 10948
rect 41076 10892 41086 10948
rect 50372 10836 50428 11116
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 30146 10780 30156 10836
rect 30212 10780 30828 10836
rect 30884 10780 30894 10836
rect 35858 10780 35868 10836
rect 35924 10780 37324 10836
rect 37380 10780 37390 10836
rect 40450 10780 40460 10836
rect 40516 10780 41356 10836
rect 41412 10780 43708 10836
rect 43764 10780 43774 10836
rect 49634 10780 49644 10836
rect 49700 10780 50428 10836
rect 12898 10668 12908 10724
rect 12964 10668 13916 10724
rect 13972 10668 14924 10724
rect 14980 10668 14990 10724
rect 23426 10668 23436 10724
rect 23492 10668 24220 10724
rect 24276 10668 25228 10724
rect 25284 10668 25294 10724
rect 31154 10668 31164 10724
rect 31220 10668 35756 10724
rect 35812 10668 35822 10724
rect 36194 10668 36204 10724
rect 36260 10668 36764 10724
rect 36820 10668 38780 10724
rect 38836 10668 39564 10724
rect 39620 10668 39630 10724
rect 42018 10668 42028 10724
rect 42084 10668 42812 10724
rect 42868 10668 42878 10724
rect 23772 10612 23828 10668
rect 42028 10612 42084 10668
rect 7074 10556 7084 10612
rect 7140 10556 10668 10612
rect 10724 10556 11116 10612
rect 11172 10556 11182 10612
rect 15250 10556 15260 10612
rect 15316 10556 16828 10612
rect 16884 10556 17500 10612
rect 17556 10556 17566 10612
rect 23762 10556 23772 10612
rect 23828 10556 23838 10612
rect 29922 10556 29932 10612
rect 29988 10556 41468 10612
rect 41524 10556 42084 10612
rect 42242 10556 42252 10612
rect 42308 10556 43820 10612
rect 43876 10556 45052 10612
rect 45108 10556 45118 10612
rect 45378 10556 45388 10612
rect 45444 10556 47964 10612
rect 48020 10556 49420 10612
rect 49476 10556 49486 10612
rect 4274 10444 4284 10500
rect 4340 10444 6188 10500
rect 6244 10444 6254 10500
rect 12450 10444 12460 10500
rect 12516 10444 13468 10500
rect 13524 10444 13534 10500
rect 33506 10444 33516 10500
rect 33572 10444 35980 10500
rect 36036 10444 36046 10500
rect 39106 10444 39116 10500
rect 39172 10444 39452 10500
rect 39508 10444 41916 10500
rect 41972 10444 41982 10500
rect 2146 10332 2156 10388
rect 2212 10332 5628 10388
rect 5684 10332 5694 10388
rect 6514 10332 6524 10388
rect 6580 10332 7420 10388
rect 7476 10332 7486 10388
rect 33394 10332 33404 10388
rect 33460 10332 35644 10388
rect 35700 10332 35710 10388
rect 26226 10220 26236 10276
rect 26292 10220 27132 10276
rect 27188 10220 27198 10276
rect 46358 10220 46396 10276
rect 46452 10220 46462 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 26002 10108 26012 10164
rect 26068 10108 29484 10164
rect 29540 10108 29550 10164
rect 36194 10108 36204 10164
rect 36260 10108 37772 10164
rect 37828 10108 37838 10164
rect 39666 10108 39676 10164
rect 39732 10108 40908 10164
rect 40964 10108 42364 10164
rect 42420 10108 42430 10164
rect 46274 10108 46284 10164
rect 46340 10108 49196 10164
rect 49252 10108 49262 10164
rect 42364 10052 42420 10108
rect 11106 9996 11116 10052
rect 11172 9996 12348 10052
rect 12404 9996 13300 10052
rect 39218 9996 39228 10052
rect 39284 9996 41132 10052
rect 41188 9996 41198 10052
rect 42364 9996 47404 10052
rect 47460 9996 47470 10052
rect 13244 9940 13300 9996
rect 11554 9884 11564 9940
rect 11620 9884 12684 9940
rect 12740 9884 12750 9940
rect 13234 9884 13244 9940
rect 13300 9884 13916 9940
rect 13972 9884 15148 9940
rect 15204 9884 15214 9940
rect 11778 9772 11788 9828
rect 11844 9772 12908 9828
rect 12964 9772 14476 9828
rect 14532 9772 15372 9828
rect 15428 9772 15438 9828
rect 16146 9772 16156 9828
rect 16212 9772 16222 9828
rect 27122 9772 27132 9828
rect 27188 9772 29148 9828
rect 29204 9772 38668 9828
rect 38724 9772 38734 9828
rect 12674 9660 12684 9716
rect 12740 9660 13580 9716
rect 13636 9660 14700 9716
rect 14756 9660 14766 9716
rect 16156 9604 16212 9772
rect 39228 9716 39284 9996
rect 43922 9772 43932 9828
rect 43988 9772 46396 9828
rect 46452 9772 46462 9828
rect 47842 9772 47852 9828
rect 47908 9772 49756 9828
rect 49812 9772 49822 9828
rect 32162 9660 32172 9716
rect 32228 9660 39284 9716
rect 45938 9660 45948 9716
rect 46004 9660 46172 9716
rect 46228 9660 48076 9716
rect 48132 9660 49084 9716
rect 49140 9660 49150 9716
rect 49858 9660 49868 9716
rect 49924 9660 50540 9716
rect 50596 9660 52780 9716
rect 52836 9660 52846 9716
rect 8082 9548 8092 9604
rect 8148 9548 11004 9604
rect 11060 9548 11070 9604
rect 11218 9548 11228 9604
rect 11284 9548 12124 9604
rect 12180 9548 12190 9604
rect 14242 9548 14252 9604
rect 14308 9548 16716 9604
rect 16772 9548 16782 9604
rect 35522 9548 35532 9604
rect 35588 9548 35980 9604
rect 36036 9548 36046 9604
rect 42690 9548 42700 9604
rect 42756 9548 43596 9604
rect 43652 9548 50092 9604
rect 50148 9548 50158 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 7410 9212 7420 9268
rect 7476 9212 21756 9268
rect 21812 9212 21822 9268
rect 35634 9212 35644 9268
rect 35700 9212 36428 9268
rect 36484 9212 36494 9268
rect 36866 9212 36876 9268
rect 36932 9212 38332 9268
rect 38388 9212 38398 9268
rect 43810 9212 43820 9268
rect 43876 9212 48300 9268
rect 48356 9212 48366 9268
rect 19618 9100 19628 9156
rect 19684 9100 23436 9156
rect 23492 9100 23502 9156
rect 31938 9100 31948 9156
rect 32004 9100 33068 9156
rect 33124 9100 33628 9156
rect 33684 9100 33694 9156
rect 35858 9100 35868 9156
rect 35924 9100 38108 9156
rect 38164 9100 38174 9156
rect 42466 8988 42476 9044
rect 42532 8988 45388 9044
rect 45444 8988 45454 9044
rect 49746 8988 49756 9044
rect 49812 8988 52220 9044
rect 52276 8988 52286 9044
rect 6066 8876 6076 8932
rect 6132 8876 9660 8932
rect 9716 8876 9726 8932
rect 31714 8764 31724 8820
rect 31780 8764 33068 8820
rect 33124 8764 33134 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 54200 8596 55000 8624
rect 20850 8540 20860 8596
rect 20916 8540 25340 8596
rect 25396 8540 25406 8596
rect 38322 8540 38332 8596
rect 38388 8540 38892 8596
rect 38948 8540 38958 8596
rect 53218 8540 53228 8596
rect 53284 8540 55000 8596
rect 54200 8512 55000 8540
rect 42130 8428 42140 8484
rect 42196 8428 42812 8484
rect 42868 8428 47292 8484
rect 47348 8428 47358 8484
rect 21746 8316 21756 8372
rect 21812 8316 26236 8372
rect 26292 8316 27244 8372
rect 27300 8316 29036 8372
rect 29092 8316 29102 8372
rect 35410 8316 35420 8372
rect 35476 8316 35756 8372
rect 35812 8316 36316 8372
rect 36372 8316 43148 8372
rect 43204 8316 44044 8372
rect 44100 8316 44110 8372
rect 5394 8204 5404 8260
rect 5460 8204 7420 8260
rect 7476 8204 8428 8260
rect 8484 8204 8494 8260
rect 20626 8204 20636 8260
rect 20692 8204 22988 8260
rect 23044 8204 23054 8260
rect 35634 8204 35644 8260
rect 35700 8204 36596 8260
rect 42914 8204 42924 8260
rect 42980 8204 43820 8260
rect 43876 8204 43886 8260
rect 46498 8204 46508 8260
rect 46564 8204 47180 8260
rect 47236 8204 48188 8260
rect 48244 8204 48254 8260
rect 36540 8148 36596 8204
rect 23202 8092 23212 8148
rect 23268 8092 23548 8148
rect 23604 8092 24556 8148
rect 24612 8092 24622 8148
rect 25442 8092 25452 8148
rect 25508 8092 26012 8148
rect 26068 8092 31388 8148
rect 31444 8092 31454 8148
rect 34962 8092 34972 8148
rect 35028 8092 35756 8148
rect 35812 8092 35822 8148
rect 36530 8092 36540 8148
rect 36596 8092 36988 8148
rect 37044 8092 37054 8148
rect 19506 7980 19516 8036
rect 19572 7980 20300 8036
rect 20356 7980 20366 8036
rect 22642 7980 22652 8036
rect 22708 7980 23100 8036
rect 23156 7980 24780 8036
rect 24836 7980 24846 8036
rect 26338 7980 26348 8036
rect 26404 7980 28700 8036
rect 28756 7980 28766 8036
rect 40786 7980 40796 8036
rect 40852 7980 42588 8036
rect 42644 7980 42654 8036
rect 39218 7868 39228 7924
rect 39284 7868 41244 7924
rect 41300 7868 41310 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 23314 7756 23324 7812
rect 23380 7756 25004 7812
rect 25060 7756 25900 7812
rect 25956 7756 25966 7812
rect 22530 7644 22540 7700
rect 22596 7644 23100 7700
rect 23156 7644 23166 7700
rect 31154 7644 31164 7700
rect 31220 7644 31836 7700
rect 31892 7644 34188 7700
rect 34244 7644 34254 7700
rect 38770 7644 38780 7700
rect 38836 7644 39004 7700
rect 39060 7644 39070 7700
rect 41458 7644 41468 7700
rect 41524 7644 42140 7700
rect 42196 7644 42206 7700
rect 45378 7644 45388 7700
rect 45444 7644 46732 7700
rect 46788 7644 46798 7700
rect 18498 7532 18508 7588
rect 18564 7532 19180 7588
rect 19236 7532 19246 7588
rect 22306 7532 22316 7588
rect 22372 7532 23436 7588
rect 23492 7532 23502 7588
rect 23762 7532 23772 7588
rect 23828 7532 36092 7588
rect 36148 7532 37884 7588
rect 37940 7532 38668 7588
rect 38724 7532 38734 7588
rect 47730 7532 47740 7588
rect 47796 7532 48300 7588
rect 48356 7532 50204 7588
rect 50260 7532 50428 7588
rect 50484 7532 52332 7588
rect 52388 7532 52398 7588
rect 8418 7420 8428 7476
rect 8484 7420 10220 7476
rect 10276 7420 10668 7476
rect 10724 7420 10734 7476
rect 18722 7420 18732 7476
rect 18788 7420 23212 7476
rect 23268 7420 23278 7476
rect 26226 7420 26236 7476
rect 26292 7420 26302 7476
rect 36978 7420 36988 7476
rect 37044 7420 37996 7476
rect 38052 7420 38062 7476
rect 46834 7420 46844 7476
rect 46900 7420 48524 7476
rect 48580 7420 48590 7476
rect 26236 7364 26292 7420
rect 8194 7308 8204 7364
rect 8260 7308 8540 7364
rect 8596 7308 8606 7364
rect 13570 7308 13580 7364
rect 13636 7308 14588 7364
rect 14644 7308 16268 7364
rect 16324 7308 17052 7364
rect 17108 7308 17948 7364
rect 18004 7308 19292 7364
rect 19348 7308 19358 7364
rect 26236 7308 26908 7364
rect 27010 7308 27020 7364
rect 27076 7308 29484 7364
rect 29540 7308 30828 7364
rect 30884 7308 31164 7364
rect 31220 7308 31230 7364
rect 32620 7308 40684 7364
rect 40740 7308 40750 7364
rect 17714 7196 17724 7252
rect 17780 7196 18396 7252
rect 18452 7196 18462 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 26852 7028 26908 7308
rect 32620 7252 32676 7308
rect 30930 7196 30940 7252
rect 30996 7196 32676 7252
rect 38612 7196 41020 7252
rect 41076 7196 41086 7252
rect 41794 7196 41804 7252
rect 41860 7196 43036 7252
rect 43092 7196 43102 7252
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 15092 6972 25452 7028
rect 25508 6972 25518 7028
rect 26852 6972 27020 7028
rect 27076 6972 31052 7028
rect 31108 6972 31118 7028
rect 15092 6916 15148 6972
rect 38612 6916 38668 7196
rect 48402 6972 48412 7028
rect 48468 6972 49196 7028
rect 49252 6972 49262 7028
rect 3602 6860 3612 6916
rect 3668 6860 15148 6916
rect 19842 6860 19852 6916
rect 19908 6860 22316 6916
rect 22372 6860 22382 6916
rect 31378 6860 31388 6916
rect 31444 6860 32844 6916
rect 32900 6860 38668 6916
rect 42466 6860 42476 6916
rect 42532 6860 43820 6916
rect 43876 6860 47684 6916
rect 47628 6804 47684 6860
rect 10658 6748 10668 6804
rect 10724 6748 12404 6804
rect 14802 6748 14812 6804
rect 14868 6748 16380 6804
rect 16436 6748 16446 6804
rect 22194 6748 22204 6804
rect 22260 6748 22988 6804
rect 23044 6748 23884 6804
rect 23940 6748 23950 6804
rect 43362 6748 43372 6804
rect 43428 6748 45108 6804
rect 12348 6692 12404 6748
rect 45052 6692 45108 6748
rect 47628 6748 49980 6804
rect 50036 6748 50046 6804
rect 47628 6692 47684 6748
rect 8978 6636 8988 6692
rect 9044 6636 9884 6692
rect 9940 6636 9950 6692
rect 12338 6636 12348 6692
rect 12404 6636 13468 6692
rect 13524 6636 13534 6692
rect 38322 6636 38332 6692
rect 38388 6636 39116 6692
rect 39172 6636 39182 6692
rect 43586 6636 43596 6692
rect 43652 6636 44828 6692
rect 44884 6636 44894 6692
rect 45052 6636 46004 6692
rect 46722 6636 46732 6692
rect 46788 6636 47404 6692
rect 47460 6636 47470 6692
rect 47618 6636 47628 6692
rect 47684 6636 47694 6692
rect 48066 6636 48076 6692
rect 48132 6636 48636 6692
rect 48692 6636 48702 6692
rect 51538 6636 51548 6692
rect 51604 6636 52668 6692
rect 52724 6636 52734 6692
rect 45948 6580 46004 6636
rect 44258 6524 44268 6580
rect 44324 6524 45724 6580
rect 45780 6524 45790 6580
rect 45948 6524 47180 6580
rect 47236 6524 49532 6580
rect 49588 6524 49598 6580
rect 9090 6412 9100 6468
rect 9156 6412 10556 6468
rect 10612 6412 10622 6468
rect 24210 6412 24220 6468
rect 24276 6412 27804 6468
rect 27860 6412 30380 6468
rect 30436 6412 31052 6468
rect 31108 6412 31118 6468
rect 44034 6412 44044 6468
rect 44100 6412 46396 6468
rect 46452 6412 47852 6468
rect 47908 6412 50204 6468
rect 50260 6412 50270 6468
rect 52210 6412 52220 6468
rect 52276 6412 53228 6468
rect 53284 6412 53294 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 22978 6076 22988 6132
rect 23044 6076 23660 6132
rect 23716 6076 24220 6132
rect 24276 6076 24286 6132
rect 24434 6076 24444 6132
rect 24500 6076 26684 6132
rect 26740 6076 27468 6132
rect 27524 6076 27534 6132
rect 24444 6020 24500 6076
rect 22530 5964 22540 6020
rect 22596 5964 22876 6020
rect 22932 5964 24500 6020
rect 54200 5908 55000 5936
rect 24546 5852 24556 5908
rect 24612 5852 27244 5908
rect 27300 5852 27692 5908
rect 27748 5852 27758 5908
rect 53330 5852 53340 5908
rect 53396 5852 55000 5908
rect 54200 5824 55000 5852
rect 19506 5740 19516 5796
rect 19572 5740 22428 5796
rect 22484 5740 22494 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 10546 5180 10556 5236
rect 10612 5180 11900 5236
rect 11956 5180 18396 5236
rect 18452 5180 18462 5236
rect 18834 5180 18844 5236
rect 18900 5180 22652 5236
rect 22708 5180 22718 5236
rect 23538 5180 23548 5236
rect 23604 5180 33404 5236
rect 33460 5180 34076 5236
rect 34132 5180 34142 5236
rect 39218 5180 39228 5236
rect 39284 5180 40908 5236
rect 40964 5180 40974 5236
rect 44370 5180 44380 5236
rect 44436 5180 44940 5236
rect 44996 5180 45006 5236
rect 16706 5068 16716 5124
rect 16772 5068 19180 5124
rect 19236 5068 19246 5124
rect 21634 5068 21644 5124
rect 21700 5068 22428 5124
rect 22484 5068 22494 5124
rect 25330 5068 25340 5124
rect 25396 5068 25788 5124
rect 25844 5068 26908 5124
rect 26964 5068 27804 5124
rect 27860 5068 28476 5124
rect 28532 5068 31276 5124
rect 31332 5068 31342 5124
rect 46722 5068 46732 5124
rect 46788 5068 48860 5124
rect 48916 5068 49980 5124
rect 50036 5068 50046 5124
rect 33954 4956 33964 5012
rect 34020 4956 35420 5012
rect 35476 4956 37324 5012
rect 37380 4956 37996 5012
rect 38052 4956 38668 5012
rect 45154 4956 45164 5012
rect 45220 4956 52668 5012
rect 52724 4956 52734 5012
rect 19282 4844 19292 4900
rect 19348 4844 21420 4900
rect 21476 4844 21486 4900
rect 28242 4844 28252 4900
rect 28308 4844 29932 4900
rect 29988 4844 29998 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 38612 4676 38668 4956
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 38612 4620 38836 4676
rect 14354 4508 14364 4564
rect 14420 4508 14924 4564
rect 14980 4508 26908 4564
rect 26852 4228 26908 4508
rect 38780 4340 38836 4620
rect 43698 4508 43708 4564
rect 43764 4508 44492 4564
rect 44548 4508 44558 4564
rect 49970 4396 49980 4452
rect 50036 4396 51100 4452
rect 51156 4396 51166 4452
rect 38770 4284 38780 4340
rect 38836 4284 41244 4340
rect 41300 4284 41310 4340
rect 26852 4172 42028 4228
rect 42084 4172 44044 4228
rect 44100 4172 44110 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 50642 3836 50652 3892
rect 50708 3836 53228 3892
rect 53284 3836 53294 3892
rect 18386 3612 18396 3668
rect 18452 3612 32900 3668
rect 34066 3612 34076 3668
rect 34132 3612 36988 3668
rect 37044 3612 37054 3668
rect 41346 3612 41356 3668
rect 41412 3612 42028 3668
rect 42084 3612 43708 3668
rect 43764 3612 43774 3668
rect 49634 3612 49644 3668
rect 49700 3612 51996 3668
rect 52052 3612 52062 3668
rect 32844 3556 32900 3612
rect 24658 3500 24668 3556
rect 24724 3500 30604 3556
rect 30660 3500 30670 3556
rect 32844 3500 35532 3556
rect 35588 3500 35980 3556
rect 36036 3500 36046 3556
rect 7186 3388 7196 3444
rect 7252 3388 10108 3444
rect 10164 3388 10174 3444
rect 11890 3388 11900 3444
rect 11956 3388 12460 3444
rect 12516 3388 23548 3444
rect 23604 3388 23614 3444
rect 38546 3388 38556 3444
rect 38612 3388 39340 3444
rect 39396 3388 39788 3444
rect 39844 3388 39854 3444
rect 43026 3388 43036 3444
rect 43092 3388 44156 3444
rect 44212 3388 44222 3444
rect 46386 3388 46396 3444
rect 46452 3388 47404 3444
rect 47460 3388 47470 3444
rect 16146 3276 16156 3332
rect 16212 3276 16940 3332
rect 16996 3276 17006 3332
rect 54200 3220 55000 3248
rect 52434 3164 52444 3220
rect 52500 3164 53228 3220
rect 53284 3164 55000 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 54200 3136 55000 3164
<< via3 >>
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 21868 50428 21924 50484
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 23548 49756 23604 49812
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 23660 49084 23716 49140
rect 23548 48636 23604 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 23660 48188 23716 48244
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 21868 47292 21924 47348
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 26348 45612 26404 45668
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 26348 35644 26404 35700
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 40012 34860 40068 34916
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 39340 29708 39396 29764
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 30716 27132 30772 27188
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 40012 26572 40068 26628
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 30716 24892 30772 24948
rect 39340 24556 39396 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 24556 21644 24612 21700
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 44268 20412 44324 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 40236 20188 40292 20244
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 44268 19404 44324 19460
rect 23996 19180 24052 19236
rect 46396 18956 46452 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 46284 17164 46340 17220
rect 24556 17052 24612 17108
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 46284 14476 46340 14532
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 46396 13692 46452 13748
rect 40236 13356 40292 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 23996 12012 24052 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 46396 10220 46452 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 46396 3388 46452 3444
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 50988 4768 51804
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 51772 20128 51804
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 35168 50988 35488 51804
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 21868 50484 21924 50494
rect 21868 47348 21924 50428
rect 23548 49812 23604 49822
rect 23548 48692 23604 49756
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 23548 48626 23604 48636
rect 23660 49140 23716 49150
rect 23660 48244 23716 49084
rect 23660 48178 23716 48188
rect 21868 47282 21924 47292
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 26348 45668 26404 45678
rect 26348 35700 26404 45612
rect 26348 35634 26404 35644
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 50528 51772 50848 51804
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 40012 34916 40068 34926
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 30716 27188 30772 27198
rect 30716 24948 30772 27132
rect 30716 24882 30772 24892
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 24332 35488 25844
rect 39340 29764 39396 29774
rect 39340 24612 39396 29708
rect 40012 26628 40068 34860
rect 40012 26562 40068 26572
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 39340 24546 39396 24556
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 24556 21700 24612 21710
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 23996 19236 24052 19246
rect 23996 12068 24052 19180
rect 24556 17108 24612 21644
rect 24556 17042 24612 17052
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 44268 20468 44324 20478
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 23996 12002 24052 12012
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 40236 20244 40292 20254
rect 40236 13412 40292 20188
rect 44268 19460 44324 20412
rect 44268 19394 44324 19404
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 46396 19012 46452 19022
rect 46284 17220 46340 17230
rect 46284 14532 46340 17164
rect 46284 14466 46340 14476
rect 46396 13748 46452 18956
rect 46396 13682 46452 13692
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 40236 13346 40292 13356
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 46396 10276 46452 10286
rect 46396 3444 46452 10220
rect 46396 3378 46452 3388
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0827_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0828_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19152 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0829_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0830_
timestamp 1698175906
transform -1 0 50064 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0831_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40096 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0832_
timestamp 1698175906
transform 1 0 38864 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0833_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0834_
timestamp 1698175906
transform -1 0 32928 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0835_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38752 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _0836_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39200 0 1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0837_
timestamp 1698175906
transform 1 0 41216 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0838_
timestamp 1698175906
transform 1 0 33824 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0839_
timestamp 1698175906
transform 1 0 36176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0840_
timestamp 1698175906
transform 1 0 37408 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0841_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0842_
timestamp 1698175906
transform -1 0 40432 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0843_
timestamp 1698175906
transform 1 0 35840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0844_
timestamp 1698175906
transform 1 0 33264 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0845_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 34496 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0846_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39872 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0847_
timestamp 1698175906
transform 1 0 36624 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0848_
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0849_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37968 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0850_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37968 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0851_
timestamp 1698175906
transform 1 0 40544 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0852_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46144 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0853_
timestamp 1698175906
transform 1 0 49168 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0854_
timestamp 1698175906
transform -1 0 42784 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0855_
timestamp 1698175906
transform -1 0 42560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0856_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40544 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0857_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 42672 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0858_
timestamp 1698175906
transform -1 0 44352 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0859_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39424 0 1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0860_
timestamp 1698175906
transform 1 0 38752 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0861_
timestamp 1698175906
transform 1 0 46256 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0862_
timestamp 1698175906
transform -1 0 47152 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0863_
timestamp 1698175906
transform -1 0 44352 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0864_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44352 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0865_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 45808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0866_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44800 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0867_
timestamp 1698175906
transform 1 0 29904 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0868_
timestamp 1698175906
transform 1 0 41328 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0869_
timestamp 1698175906
transform 1 0 46032 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0870_
timestamp 1698175906
transform -1 0 47824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0871_
timestamp 1698175906
transform -1 0 47376 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0872_
timestamp 1698175906
transform 1 0 47264 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0873_
timestamp 1698175906
transform -1 0 49280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0874_
timestamp 1698175906
transform 1 0 49280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0875_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 47152 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0876_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 46256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0877_
timestamp 1698175906
transform 1 0 46480 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0878_
timestamp 1698175906
transform -1 0 41664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0879_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 41104 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0880_
timestamp 1698175906
transform -1 0 43456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0881_
timestamp 1698175906
transform -1 0 50960 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0882_
timestamp 1698175906
transform 1 0 46032 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0883_
timestamp 1698175906
transform 1 0 49056 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0884_
timestamp 1698175906
transform 1 0 49392 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0885_
timestamp 1698175906
transform 1 0 49504 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0886_
timestamp 1698175906
transform 1 0 48496 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0887_
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698175906
transform 1 0 51744 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0889_
timestamp 1698175906
transform 1 0 50400 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0891_
timestamp 1698175906
transform 1 0 51072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0892_
timestamp 1698175906
transform 1 0 51968 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0893_
timestamp 1698175906
transform 1 0 49392 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0894_
timestamp 1698175906
transform 1 0 51520 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0895_
timestamp 1698175906
transform 1 0 50960 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0896_
timestamp 1698175906
transform 1 0 52192 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0897_
timestamp 1698175906
transform 1 0 51296 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0898_
timestamp 1698175906
transform -1 0 51296 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0899_
timestamp 1698175906
transform -1 0 46032 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0900_
timestamp 1698175906
transform 1 0 43344 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0901_
timestamp 1698175906
transform -1 0 50624 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0902_
timestamp 1698175906
transform 1 0 49504 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0903_
timestamp 1698175906
transform 1 0 49728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0904_
timestamp 1698175906
transform -1 0 51744 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0905_
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0906_
timestamp 1698175906
transform 1 0 50400 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0907_
timestamp 1698175906
transform 1 0 49616 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0908_
timestamp 1698175906
transform -1 0 51856 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0909_
timestamp 1698175906
transform 1 0 51296 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0910_
timestamp 1698175906
transform 1 0 51408 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0911_
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0912_
timestamp 1698175906
transform 1 0 48944 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0913_
timestamp 1698175906
transform 1 0 49168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0914_
timestamp 1698175906
transform -1 0 50960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0915_
timestamp 1698175906
transform -1 0 47152 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0916_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 52976 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0917_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 48608 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0918_
timestamp 1698175906
transform -1 0 42560 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0919_
timestamp 1698175906
transform -1 0 44240 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0920_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 46256 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0921_
timestamp 1698175906
transform 1 0 42000 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0922_
timestamp 1698175906
transform 1 0 49056 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0923_
timestamp 1698175906
transform 1 0 50512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0924_
timestamp 1698175906
transform -1 0 52864 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0925_
timestamp 1698175906
transform -1 0 50736 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0926_
timestamp 1698175906
transform -1 0 50624 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0927_
timestamp 1698175906
transform -1 0 44240 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0928_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 49392 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0929_
timestamp 1698175906
transform 1 0 50624 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0930_
timestamp 1698175906
transform -1 0 49504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0931_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 48160 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0932_
timestamp 1698175906
transform 1 0 48272 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0933_
timestamp 1698175906
transform -1 0 47040 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0934_
timestamp 1698175906
transform 1 0 47040 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0935_
timestamp 1698175906
transform -1 0 47824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0936_
timestamp 1698175906
transform -1 0 46816 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0937_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46144 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0938_
timestamp 1698175906
transform 1 0 43232 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0939_
timestamp 1698175906
transform -1 0 45136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0940_
timestamp 1698175906
transform 1 0 31360 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0941_
timestamp 1698175906
transform 1 0 45136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0942_
timestamp 1698175906
transform -1 0 42336 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0943_
timestamp 1698175906
transform -1 0 50624 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1698175906
transform 1 0 42000 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0945_
timestamp 1698175906
transform -1 0 46256 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0946_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46144 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0947_
timestamp 1698175906
transform -1 0 45248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0948_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 45024 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0949_
timestamp 1698175906
transform -1 0 20944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0950_
timestamp 1698175906
transform 1 0 24640 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0951_
timestamp 1698175906
transform -1 0 29680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0952_
timestamp 1698175906
transform -1 0 26432 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0953_
timestamp 1698175906
transform -1 0 30016 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0954_
timestamp 1698175906
transform -1 0 29568 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0955_
timestamp 1698175906
transform 1 0 26768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0956_
timestamp 1698175906
transform -1 0 34160 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0957_
timestamp 1698175906
transform -1 0 41664 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0958_
timestamp 1698175906
transform -1 0 39872 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0959_
timestamp 1698175906
transform -1 0 36960 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0960_
timestamp 1698175906
transform -1 0 33600 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0961_
timestamp 1698175906
transform -1 0 32368 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0962_
timestamp 1698175906
transform -1 0 34832 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0963_
timestamp 1698175906
transform 1 0 37744 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698175906
transform 1 0 38528 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0965_
timestamp 1698175906
transform 1 0 31696 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0966_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32032 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0967_
timestamp 1698175906
transform -1 0 44464 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0968_
timestamp 1698175906
transform -1 0 32032 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0969_
timestamp 1698175906
transform 1 0 31584 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0970_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 34720 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0971_
timestamp 1698175906
transform 1 0 35616 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0972_
timestamp 1698175906
transform 1 0 26320 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0973_
timestamp 1698175906
transform -1 0 32480 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0974_
timestamp 1698175906
transform 1 0 38528 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0975_
timestamp 1698175906
transform 1 0 35504 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0976_
timestamp 1698175906
transform 1 0 39536 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0977_
timestamp 1698175906
transform 1 0 41776 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0978_
timestamp 1698175906
transform 1 0 45136 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0979_
timestamp 1698175906
transform 1 0 35280 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0980_
timestamp 1698175906
transform 1 0 38416 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0981_
timestamp 1698175906
transform 1 0 40320 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0982_
timestamp 1698175906
transform 1 0 42112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0983_
timestamp 1698175906
transform -1 0 37520 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0984_
timestamp 1698175906
transform -1 0 38528 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0985_
timestamp 1698175906
transform -1 0 36400 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0986_
timestamp 1698175906
transform -1 0 36064 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0987_
timestamp 1698175906
transform -1 0 36064 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0988_
timestamp 1698175906
transform -1 0 35168 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0989_
timestamp 1698175906
transform 1 0 36064 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0990_
timestamp 1698175906
transform 1 0 37968 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0991_
timestamp 1698175906
transform -1 0 39424 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0992_
timestamp 1698175906
transform -1 0 38528 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0993_
timestamp 1698175906
transform -1 0 20720 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0994_
timestamp 1698175906
transform 1 0 23296 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0995_
timestamp 1698175906
transform -1 0 37072 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0996_
timestamp 1698175906
transform 1 0 38976 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0997_
timestamp 1698175906
transform 1 0 38864 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0998_
timestamp 1698175906
transform -1 0 39424 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0999_
timestamp 1698175906
transform 1 0 39648 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1000_
timestamp 1698175906
transform -1 0 30912 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1001_
timestamp 1698175906
transform 1 0 30912 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1002_
timestamp 1698175906
transform -1 0 42000 0 -1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1003_
timestamp 1698175906
transform -1 0 43568 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1004_
timestamp 1698175906
transform 1 0 40656 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1005_
timestamp 1698175906
transform 1 0 25984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1006_
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1007_
timestamp 1698175906
transform 1 0 26432 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1008_
timestamp 1698175906
transform -1 0 26880 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698175906
transform -1 0 29344 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1010_
timestamp 1698175906
transform 1 0 24192 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1011_
timestamp 1698175906
transform 1 0 25872 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1012_
timestamp 1698175906
transform -1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1013_
timestamp 1698175906
transform -1 0 24864 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1014_
timestamp 1698175906
transform -1 0 24528 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1015_
timestamp 1698175906
transform -1 0 24304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1016_
timestamp 1698175906
transform -1 0 25760 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1017_
timestamp 1698175906
transform 1 0 23296 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698175906
transform -1 0 25984 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1019_
timestamp 1698175906
transform -1 0 23632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1020_
timestamp 1698175906
transform -1 0 25872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1021_
timestamp 1698175906
transform -1 0 23520 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1022_
timestamp 1698175906
transform -1 0 24528 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1023_
timestamp 1698175906
transform -1 0 23744 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1024_
timestamp 1698175906
transform -1 0 23856 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1025_
timestamp 1698175906
transform -1 0 24192 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1026_
timestamp 1698175906
transform -1 0 23968 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1027_
timestamp 1698175906
transform -1 0 24416 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1028_
timestamp 1698175906
transform -1 0 24304 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1029_
timestamp 1698175906
transform 1 0 23632 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1030_
timestamp 1698175906
transform 1 0 26992 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1031_
timestamp 1698175906
transform 1 0 26656 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1032_
timestamp 1698175906
transform -1 0 30688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1033_
timestamp 1698175906
transform 1 0 25200 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1034_
timestamp 1698175906
transform 1 0 26096 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1035_
timestamp 1698175906
transform 1 0 27328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1036_
timestamp 1698175906
transform -1 0 36288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1037_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32256 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1038_
timestamp 1698175906
transform -1 0 32480 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1039_
timestamp 1698175906
transform -1 0 44464 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1040_
timestamp 1698175906
transform -1 0 29680 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1041_
timestamp 1698175906
transform -1 0 44800 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1042_
timestamp 1698175906
transform -1 0 39872 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1043_
timestamp 1698175906
transform -1 0 37408 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1044_
timestamp 1698175906
transform -1 0 31024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1045_
timestamp 1698175906
transform -1 0 32032 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1046_
timestamp 1698175906
transform 1 0 35392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698175906
transform -1 0 35392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1048_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30800 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1049_
timestamp 1698175906
transform -1 0 31248 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1050_
timestamp 1698175906
transform 1 0 30352 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1051_
timestamp 1698175906
transform -1 0 34720 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1052_
timestamp 1698175906
transform -1 0 45248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1053_
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1054_
timestamp 1698175906
transform -1 0 34720 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1055_
timestamp 1698175906
transform -1 0 31584 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1056_
timestamp 1698175906
transform 1 0 31472 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1057_
timestamp 1698175906
transform -1 0 31472 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1058_
timestamp 1698175906
transform -1 0 45360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1059_
timestamp 1698175906
transform -1 0 31584 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1060_
timestamp 1698175906
transform 1 0 30576 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1061_
timestamp 1698175906
transform 1 0 31136 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1062_
timestamp 1698175906
transform 1 0 34384 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1063_
timestamp 1698175906
transform -1 0 43344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1064_
timestamp 1698175906
transform 1 0 34048 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1065_
timestamp 1698175906
transform 1 0 32928 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1066_
timestamp 1698175906
transform 1 0 33264 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1067_
timestamp 1698175906
transform 1 0 33936 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1068_
timestamp 1698175906
transform -1 0 49504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1069_
timestamp 1698175906
transform 1 0 33488 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1070_
timestamp 1698175906
transform 1 0 33152 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1071_
timestamp 1698175906
transform 1 0 33600 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698175906
transform -1 0 45360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1073_
timestamp 1698175906
transform 1 0 34720 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1074_
timestamp 1698175906
transform 1 0 33824 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1075_
timestamp 1698175906
transform 1 0 35392 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1076_
timestamp 1698175906
transform -1 0 49840 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1077_
timestamp 1698175906
transform 1 0 34720 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1078_
timestamp 1698175906
transform 1 0 33824 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1079_
timestamp 1698175906
transform 1 0 34608 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 47824 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1081_
timestamp 1698175906
transform 1 0 49504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1082_
timestamp 1698175906
transform 1 0 44016 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1083_
timestamp 1698175906
transform 1 0 48608 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1084_
timestamp 1698175906
transform -1 0 39200 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1085_
timestamp 1698175906
transform -1 0 43792 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1086_
timestamp 1698175906
transform 1 0 42000 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1087_
timestamp 1698175906
transform 1 0 42560 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1088_
timestamp 1698175906
transform -1 0 39536 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1089_
timestamp 1698175906
transform 1 0 43120 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1090_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 43344 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1091_
timestamp 1698175906
transform 1 0 27888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1092_
timestamp 1698175906
transform 1 0 43008 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1093_
timestamp 1698175906
transform 1 0 43456 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1094_
timestamp 1698175906
transform -1 0 46256 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1095_
timestamp 1698175906
transform 1 0 41664 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1096_
timestamp 1698175906
transform 1 0 42336 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1097_
timestamp 1698175906
transform 1 0 29232 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1098_
timestamp 1698175906
transform 1 0 41664 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1099_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 33824 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1100_
timestamp 1698175906
transform 1 0 40768 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1101_
timestamp 1698175906
transform -1 0 40544 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1102_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39648 0 -1 21952
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1103_
timestamp 1698175906
transform 1 0 44800 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1104_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 48720 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1105_
timestamp 1698175906
transform 1 0 50064 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1106_
timestamp 1698175906
transform -1 0 42336 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1107_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32704 0 -1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1108_
timestamp 1698175906
transform 1 0 38752 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1109_
timestamp 1698175906
transform -1 0 45584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1110_
timestamp 1698175906
transform 1 0 30688 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1698175906
transform 1 0 36960 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1112_
timestamp 1698175906
transform -1 0 41664 0 1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1113_
timestamp 1698175906
transform -1 0 45360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1114_
timestamp 1698175906
transform -1 0 49952 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1115_
timestamp 1698175906
transform 1 0 44912 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1116_
timestamp 1698175906
transform -1 0 33600 0 1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1117_
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1118_
timestamp 1698175906
transform 1 0 36960 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1119_
timestamp 1698175906
transform -1 0 41664 0 1 20384
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1120_
timestamp 1698175906
transform -1 0 49840 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1698175906
transform 1 0 45472 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1122_
timestamp 1698175906
transform 1 0 49280 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1123_
timestamp 1698175906
transform -1 0 42560 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1124_
timestamp 1698175906
transform -1 0 29904 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698175906
transform 1 0 27776 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1126_
timestamp 1698175906
transform -1 0 38304 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1127_
timestamp 1698175906
transform 1 0 41664 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1128_
timestamp 1698175906
transform -1 0 50512 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1129_
timestamp 1698175906
transform 1 0 50736 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1130_
timestamp 1698175906
transform 1 0 42336 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1131_
timestamp 1698175906
transform -1 0 27776 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1132_
timestamp 1698175906
transform 1 0 23408 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1133_
timestamp 1698175906
transform -1 0 40432 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1134_
timestamp 1698175906
transform -1 0 39760 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1135_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 41776 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1136_
timestamp 1698175906
transform -1 0 51408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1137_
timestamp 1698175906
transform 1 0 50736 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1138_
timestamp 1698175906
transform 1 0 30912 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1139_
timestamp 1698175906
transform 1 0 48720 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1140_
timestamp 1698175906
transform 1 0 43568 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1141_
timestamp 1698175906
transform 1 0 23072 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1142_
timestamp 1698175906
transform 1 0 38080 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1143_
timestamp 1698175906
transform 1 0 42784 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1144_
timestamp 1698175906
transform -1 0 50176 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1145_
timestamp 1698175906
transform 1 0 50512 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1146_
timestamp 1698175906
transform 1 0 44688 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1147_
timestamp 1698175906
transform 1 0 23520 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1148_
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1149_
timestamp 1698175906
transform 1 0 43568 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1150_
timestamp 1698175906
transform -1 0 50176 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1151_
timestamp 1698175906
transform 1 0 50400 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1152_
timestamp 1698175906
transform 1 0 40432 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1153_
timestamp 1698175906
transform 1 0 26656 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1154_
timestamp 1698175906
transform -1 0 39648 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1155_
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1156_
timestamp 1698175906
transform -1 0 51520 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1157_
timestamp 1698175906
transform 1 0 51520 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1158_
timestamp 1698175906
transform -1 0 34048 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1159_
timestamp 1698175906
transform 1 0 18144 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1160_
timestamp 1698175906
transform 1 0 18704 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1161_
timestamp 1698175906
transform 1 0 17360 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1162_
timestamp 1698175906
transform 1 0 17360 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1163_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1164_
timestamp 1698175906
transform 1 0 12992 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1165_
timestamp 1698175906
transform -1 0 21056 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1166_
timestamp 1698175906
transform 1 0 15680 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1167_
timestamp 1698175906
transform 1 0 14336 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1168_
timestamp 1698175906
transform 1 0 16464 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1169_
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1170_
timestamp 1698175906
transform 1 0 28112 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1171_
timestamp 1698175906
transform 1 0 27440 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1172_
timestamp 1698175906
transform 1 0 27440 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1173_
timestamp 1698175906
transform 1 0 26768 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1174_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30128 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1175_
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1176_
timestamp 1698175906
transform 1 0 21728 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1177_
timestamp 1698175906
transform 1 0 22848 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1178_
timestamp 1698175906
transform 1 0 21504 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1179_
timestamp 1698175906
transform 1 0 24192 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1180_
timestamp 1698175906
transform 1 0 28896 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1181_
timestamp 1698175906
transform 1 0 32256 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1182_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 47040 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1183_
timestamp 1698175906
transform 1 0 33376 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1184_
timestamp 1698175906
transform -1 0 39200 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1185_
timestamp 1698175906
transform 1 0 38080 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1186_
timestamp 1698175906
transform 1 0 46032 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1187_
timestamp 1698175906
transform -1 0 47040 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1188_
timestamp 1698175906
transform 1 0 48608 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1189_
timestamp 1698175906
transform 1 0 49168 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1190_
timestamp 1698175906
transform 1 0 50624 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1191_
timestamp 1698175906
transform 1 0 48720 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1192_
timestamp 1698175906
transform 1 0 48608 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1193_
timestamp 1698175906
transform -1 0 50176 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1194_
timestamp 1698175906
transform 1 0 51072 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1195_
timestamp 1698175906
transform -1 0 49056 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1196_
timestamp 1698175906
transform 1 0 47600 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1197_
timestamp 1698175906
transform -1 0 49392 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1198_
timestamp 1698175906
transform -1 0 48384 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1199_
timestamp 1698175906
transform -1 0 48944 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1200_
timestamp 1698175906
transform 1 0 46928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1201_
timestamp 1698175906
transform 1 0 47264 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1202_
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1203_
timestamp 1698175906
transform 1 0 46256 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1204_
timestamp 1698175906
transform -1 0 47712 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1205_
timestamp 1698175906
transform 1 0 46704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1206_
timestamp 1698175906
transform 1 0 47712 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1207_
timestamp 1698175906
transform 1 0 27776 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1208_
timestamp 1698175906
transform 1 0 25760 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1209_
timestamp 1698175906
transform -1 0 27104 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1210_
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1211_
timestamp 1698175906
transform 1 0 29344 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1212_
timestamp 1698175906
transform 1 0 28224 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1213_
timestamp 1698175906
transform -1 0 27888 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1214_
timestamp 1698175906
transform -1 0 27888 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1215_
timestamp 1698175906
transform -1 0 25872 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1216_
timestamp 1698175906
transform 1 0 26208 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1217_
timestamp 1698175906
transform 1 0 26880 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1218_
timestamp 1698175906
transform -1 0 26656 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1219_
timestamp 1698175906
transform 1 0 25312 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1220_
timestamp 1698175906
transform 1 0 25872 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1221_
timestamp 1698175906
transform -1 0 24640 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1222_
timestamp 1698175906
transform -1 0 22848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698175906
transform -1 0 22848 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1224_
timestamp 1698175906
transform -1 0 24864 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1225_
timestamp 1698175906
transform 1 0 21392 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1226_
timestamp 1698175906
transform -1 0 22288 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1227_
timestamp 1698175906
transform -1 0 22176 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1228_
timestamp 1698175906
transform 1 0 21728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1229_
timestamp 1698175906
transform -1 0 22736 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1230_
timestamp 1698175906
transform -1 0 22064 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1231_
timestamp 1698175906
transform 1 0 21280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1232_
timestamp 1698175906
transform -1 0 24416 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1233_
timestamp 1698175906
transform 1 0 22400 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1234_
timestamp 1698175906
transform 1 0 22960 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1235_
timestamp 1698175906
transform -1 0 38192 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1236_
timestamp 1698175906
transform 1 0 38864 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1237_
timestamp 1698175906
transform 1 0 38192 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1238_
timestamp 1698175906
transform -1 0 35168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1239_
timestamp 1698175906
transform -1 0 35168 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1240_
timestamp 1698175906
transform -1 0 37408 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1241_
timestamp 1698175906
transform -1 0 36512 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1242_
timestamp 1698175906
transform 1 0 37632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1698175906
transform -1 0 35056 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1244_
timestamp 1698175906
transform 1 0 33488 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1245_
timestamp 1698175906
transform -1 0 34608 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1246_
timestamp 1698175906
transform -1 0 32704 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1247_
timestamp 1698175906
transform -1 0 32144 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1248_
timestamp 1698175906
transform 1 0 39984 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1249_
timestamp 1698175906
transform 1 0 40544 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1698175906
transform 1 0 25648 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1251_
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1252_
timestamp 1698175906
transform 1 0 36064 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1253_
timestamp 1698175906
transform -1 0 38304 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1254_
timestamp 1698175906
transform -1 0 37744 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1255_
timestamp 1698175906
transform 1 0 39872 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1256_
timestamp 1698175906
transform 1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1257_
timestamp 1698175906
transform 1 0 39984 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1258_
timestamp 1698175906
transform 1 0 39200 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1259_
timestamp 1698175906
transform 1 0 39648 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1260_
timestamp 1698175906
transform -1 0 31696 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1261_
timestamp 1698175906
transform -1 0 24416 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1262_
timestamp 1698175906
transform -1 0 35392 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1263_
timestamp 1698175906
transform 1 0 28112 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1264_
timestamp 1698175906
transform 1 0 32928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1265_
timestamp 1698175906
transform 1 0 31696 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1266_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 34608 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1267_
timestamp 1698175906
transform 1 0 23968 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1268_
timestamp 1698175906
transform 1 0 23408 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1269_
timestamp 1698175906
transform -1 0 25760 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1270_
timestamp 1698175906
transform 1 0 26208 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1271_
timestamp 1698175906
transform 1 0 20048 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1272_
timestamp 1698175906
transform -1 0 25984 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1273_
timestamp 1698175906
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1274_
timestamp 1698175906
transform -1 0 35280 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1275_
timestamp 1698175906
transform -1 0 34720 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1698175906
transform -1 0 22960 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1277_
timestamp 1698175906
transform 1 0 24080 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1278_
timestamp 1698175906
transform 1 0 25088 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1279_
timestamp 1698175906
transform -1 0 24752 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1280_
timestamp 1698175906
transform 1 0 14224 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1281_
timestamp 1698175906
transform -1 0 21952 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1282_
timestamp 1698175906
transform -1 0 19936 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1283_
timestamp 1698175906
transform 1 0 19824 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1284_
timestamp 1698175906
transform -1 0 23744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1285_
timestamp 1698175906
transform -1 0 23072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1286_
timestamp 1698175906
transform 1 0 18928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1287_
timestamp 1698175906
transform 1 0 17584 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698175906
transform -1 0 20608 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1289_
timestamp 1698175906
transform 1 0 20720 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1290_
timestamp 1698175906
transform -1 0 21840 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1291_
timestamp 1698175906
transform -1 0 19376 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1292_
timestamp 1698175906
transform 1 0 17584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1293_
timestamp 1698175906
transform 1 0 18144 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1294_
timestamp 1698175906
transform 1 0 20272 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1295_
timestamp 1698175906
transform 1 0 21616 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1296_
timestamp 1698175906
transform -1 0 38752 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1297_
timestamp 1698175906
transform 1 0 23296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1298_
timestamp 1698175906
transform -1 0 21504 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1698175906
transform 1 0 17472 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1300_
timestamp 1698175906
transform 1 0 19488 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1301_
timestamp 1698175906
transform -1 0 26432 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1302_
timestamp 1698175906
transform 1 0 21168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1303_
timestamp 1698175906
transform -1 0 24976 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1304_
timestamp 1698175906
transform 1 0 21392 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1305_
timestamp 1698175906
transform 1 0 22288 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1306_
timestamp 1698175906
transform 1 0 27776 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1307_
timestamp 1698175906
transform -1 0 24528 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1308_
timestamp 1698175906
transform -1 0 25984 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1309_
timestamp 1698175906
transform 1 0 25760 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1310_
timestamp 1698175906
transform -1 0 23744 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1311_
timestamp 1698175906
transform -1 0 23408 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1312_
timestamp 1698175906
transform 1 0 26096 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1313_
timestamp 1698175906
transform 1 0 27216 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1314_
timestamp 1698175906
transform 1 0 25648 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1315_
timestamp 1698175906
transform 1 0 25984 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1316_
timestamp 1698175906
transform 1 0 26320 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1317_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24640 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1318_
timestamp 1698175906
transform -1 0 22848 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1319_
timestamp 1698175906
transform -1 0 29344 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1320_
timestamp 1698175906
transform -1 0 22400 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1321_
timestamp 1698175906
transform 1 0 22848 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1322_
timestamp 1698175906
transform 1 0 22960 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1323_
timestamp 1698175906
transform 1 0 22400 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1324_
timestamp 1698175906
transform 1 0 25760 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1325_
timestamp 1698175906
transform 1 0 19264 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1326_
timestamp 1698175906
transform -1 0 20832 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1327_
timestamp 1698175906
transform -1 0 21280 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1328_
timestamp 1698175906
transform 1 0 20160 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1329_
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1330_
timestamp 1698175906
transform -1 0 20272 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1331_
timestamp 1698175906
transform 1 0 17136 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698175906
transform -1 0 17808 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1333_
timestamp 1698175906
transform -1 0 16576 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1334_
timestamp 1698175906
transform 1 0 16128 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1335_
timestamp 1698175906
transform -1 0 17696 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1336_
timestamp 1698175906
transform 1 0 16576 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1337_
timestamp 1698175906
transform -1 0 16576 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1338_
timestamp 1698175906
transform 1 0 16016 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1339_
timestamp 1698175906
transform 1 0 18592 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1340_
timestamp 1698175906
transform -1 0 25312 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1341_
timestamp 1698175906
transform 1 0 10640 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14112 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1343_
timestamp 1698175906
transform -1 0 11984 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1344_
timestamp 1698175906
transform 1 0 10528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1345_
timestamp 1698175906
transform 1 0 10752 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1346_
timestamp 1698175906
transform 1 0 9856 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1347_
timestamp 1698175906
transform 1 0 9520 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1348_
timestamp 1698175906
transform 1 0 10752 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1349_
timestamp 1698175906
transform -1 0 14560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1350_
timestamp 1698175906
transform 1 0 11648 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1351_
timestamp 1698175906
transform -1 0 11200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1352_
timestamp 1698175906
transform 1 0 10640 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1353_
timestamp 1698175906
transform -1 0 13104 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1354_
timestamp 1698175906
transform 1 0 11984 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1355_
timestamp 1698175906
transform 1 0 12320 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1356_
timestamp 1698175906
transform -1 0 13664 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1357_
timestamp 1698175906
transform -1 0 11424 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1358_
timestamp 1698175906
transform -1 0 10864 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1359_
timestamp 1698175906
transform -1 0 14896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1360_
timestamp 1698175906
transform 1 0 12320 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1361_
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1362_
timestamp 1698175906
transform -1 0 20272 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1363_
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1364_
timestamp 1698175906
transform -1 0 50064 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1365_
timestamp 1698175906
transform 1 0 35392 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1366_
timestamp 1698175906
transform 1 0 37520 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1367_
timestamp 1698175906
transform -1 0 39536 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1368_
timestamp 1698175906
transform -1 0 39648 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1698175906
transform -1 0 37520 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1370_
timestamp 1698175906
transform -1 0 35280 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_
timestamp 1698175906
transform -1 0 33600 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1372_
timestamp 1698175906
transform -1 0 43008 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1373_
timestamp 1698175906
transform -1 0 35280 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1698175906
transform -1 0 34272 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1375_
timestamp 1698175906
transform -1 0 37408 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1376_
timestamp 1698175906
transform 1 0 37408 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1698175906
transform 1 0 38976 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1378_
timestamp 1698175906
transform -1 0 40432 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1379_
timestamp 1698175906
transform 1 0 40768 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1380_
timestamp 1698175906
transform -1 0 43232 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1381_
timestamp 1698175906
transform -1 0 42560 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1382_
timestamp 1698175906
transform 1 0 41328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1383_
timestamp 1698175906
transform 1 0 42224 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1384_
timestamp 1698175906
transform 1 0 42560 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1385_
timestamp 1698175906
transform 1 0 41440 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1386_
timestamp 1698175906
transform 1 0 42112 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1387_
timestamp 1698175906
transform -1 0 37296 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1388_
timestamp 1698175906
transform -1 0 37744 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1389_
timestamp 1698175906
transform 1 0 31696 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1390_
timestamp 1698175906
transform 1 0 39648 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1391_
timestamp 1698175906
transform -1 0 38752 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1392_
timestamp 1698175906
transform -1 0 29904 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1393_
timestamp 1698175906
transform -1 0 16240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1394_
timestamp 1698175906
transform 1 0 15008 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1395_
timestamp 1698175906
transform 1 0 15344 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1396_
timestamp 1698175906
transform -1 0 16688 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1397_
timestamp 1698175906
transform -1 0 16352 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1398_
timestamp 1698175906
transform -1 0 15344 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1399_
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1400_
timestamp 1698175906
transform 1 0 11536 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1401_
timestamp 1698175906
transform 1 0 12432 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1402_
timestamp 1698175906
transform 1 0 11088 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1403_
timestamp 1698175906
transform 1 0 12880 0 -1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1404_
timestamp 1698175906
transform 1 0 14896 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1405_
timestamp 1698175906
transform -1 0 8848 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1406_
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1407_
timestamp 1698175906
transform 1 0 19152 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1408_
timestamp 1698175906
transform 1 0 17136 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1409_
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1410_
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1411_
timestamp 1698175906
transform 1 0 17920 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1412_
timestamp 1698175906
transform 1 0 17696 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1413_
timestamp 1698175906
transform 1 0 17472 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1414_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1415_
timestamp 1698175906
transform -1 0 19936 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1698175906
transform -1 0 18816 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1417_
timestamp 1698175906
transform -1 0 8512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1418_
timestamp 1698175906
transform 1 0 4816 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1419_
timestamp 1698175906
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1420_
timestamp 1698175906
transform -1 0 32256 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1421_
timestamp 1698175906
transform -1 0 9408 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1422_
timestamp 1698175906
transform 1 0 7952 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1423_
timestamp 1698175906
transform -1 0 6160 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1424_
timestamp 1698175906
transform 1 0 5040 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1425_
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1426_
timestamp 1698175906
transform -1 0 7616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1427_
timestamp 1698175906
transform 1 0 10080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1428_
timestamp 1698175906
transform -1 0 10080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1429_
timestamp 1698175906
transform -1 0 9184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698175906
transform -1 0 8736 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1431_
timestamp 1698175906
transform -1 0 9184 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1432_
timestamp 1698175906
transform -1 0 2800 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1433_
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1434_
timestamp 1698175906
transform -1 0 32592 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1435_
timestamp 1698175906
transform -1 0 15232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1436_
timestamp 1698175906
transform -1 0 12880 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1437_
timestamp 1698175906
transform 1 0 6048 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1438_
timestamp 1698175906
transform 1 0 7168 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1439_
timestamp 1698175906
transform 1 0 7504 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1440_
timestamp 1698175906
transform 1 0 8176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1441_
timestamp 1698175906
transform -1 0 7504 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1442_
timestamp 1698175906
transform 1 0 3920 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1443_
timestamp 1698175906
transform 1 0 5824 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698175906
transform 1 0 9968 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1445_
timestamp 1698175906
transform -1 0 7056 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1446_
timestamp 1698175906
transform 1 0 6160 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1447_
timestamp 1698175906
transform 1 0 5488 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1448_
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1449_
timestamp 1698175906
transform 1 0 9520 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1450_
timestamp 1698175906
transform 1 0 14112 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1698175906
transform -1 0 11424 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1452_
timestamp 1698175906
transform -1 0 7168 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698175906
transform -1 0 10864 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1454_
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1455_
timestamp 1698175906
transform -1 0 11760 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1456_
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1457_
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1458_
timestamp 1698175906
transform -1 0 13104 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1459_
timestamp 1698175906
transform 1 0 10976 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1460_
timestamp 1698175906
transform 1 0 11424 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1461_
timestamp 1698175906
transform 1 0 10528 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1462_
timestamp 1698175906
transform -1 0 11984 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1463_
timestamp 1698175906
transform -1 0 15008 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698175906
transform -1 0 15904 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1465_
timestamp 1698175906
transform -1 0 13104 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1466_
timestamp 1698175906
transform -1 0 14448 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1467_
timestamp 1698175906
transform -1 0 13104 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1468_
timestamp 1698175906
transform -1 0 17024 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1469_
timestamp 1698175906
transform 1 0 13440 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1470_
timestamp 1698175906
transform -1 0 14112 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1471_
timestamp 1698175906
transform -1 0 14560 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1472_
timestamp 1698175906
transform -1 0 14672 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1473_
timestamp 1698175906
transform -1 0 19040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1474_
timestamp 1698175906
transform 1 0 14896 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1475_
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1476_
timestamp 1698175906
transform -1 0 16576 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1478_
timestamp 1698175906
transform 1 0 15456 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1479_
timestamp 1698175906
transform -1 0 21168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1480_
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698175906
transform 1 0 15568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1482_
timestamp 1698175906
transform 1 0 18144 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1483_
timestamp 1698175906
transform 1 0 17024 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1484_
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1485_
timestamp 1698175906
transform -1 0 20384 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1486_
timestamp 1698175906
transform 1 0 18144 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1487_
timestamp 1698175906
transform 1 0 17024 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1488_
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1489_
timestamp 1698175906
transform 1 0 15568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1490_
timestamp 1698175906
transform 1 0 17136 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1491_
timestamp 1698175906
transform 1 0 15904 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1492_
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1493_
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1494_
timestamp 1698175906
transform -1 0 15904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1495_
timestamp 1698175906
transform 1 0 14336 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1496_
timestamp 1698175906
transform -1 0 17136 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1497_
timestamp 1698175906
transform -1 0 14112 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1498_
timestamp 1698175906
transform 1 0 10192 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1698175906
transform -1 0 10864 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1500_
timestamp 1698175906
transform 1 0 6384 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1501_
timestamp 1698175906
transform 1 0 11312 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1502_
timestamp 1698175906
transform -1 0 12096 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1503_
timestamp 1698175906
transform -1 0 7616 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1504_
timestamp 1698175906
transform 1 0 6496 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1505_
timestamp 1698175906
transform 1 0 8512 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1506_
timestamp 1698175906
transform -1 0 11200 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1507_
timestamp 1698175906
transform 1 0 12544 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1508_
timestamp 1698175906
transform -1 0 12432 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1509_
timestamp 1698175906
transform -1 0 10304 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1510_
timestamp 1698175906
transform -1 0 10416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1511_
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1512_
timestamp 1698175906
transform -1 0 10080 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1513_
timestamp 1698175906
transform 1 0 9184 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1514_
timestamp 1698175906
transform -1 0 10304 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1515_
timestamp 1698175906
transform -1 0 10416 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1516_
timestamp 1698175906
transform -1 0 15792 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1517_
timestamp 1698175906
transform -1 0 12656 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1518_
timestamp 1698175906
transform 1 0 10192 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1519_
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1520_
timestamp 1698175906
transform 1 0 10976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1521_
timestamp 1698175906
transform 1 0 12208 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1522_
timestamp 1698175906
transform -1 0 13776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1523_
timestamp 1698175906
transform -1 0 13104 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1524_
timestamp 1698175906
transform 1 0 10752 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1525_
timestamp 1698175906
transform 1 0 11088 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1526_
timestamp 1698175906
transform 1 0 12208 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1698175906
transform -1 0 9184 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1528_
timestamp 1698175906
transform 1 0 7840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1529_
timestamp 1698175906
transform -1 0 8400 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1530_
timestamp 1698175906
transform -1 0 8176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698175906
transform -1 0 7728 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1532_
timestamp 1698175906
transform -1 0 6160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1533_
timestamp 1698175906
transform 1 0 5152 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1534_
timestamp 1698175906
transform 1 0 6272 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1535_
timestamp 1698175906
transform -1 0 9744 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1536_
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1537_
timestamp 1698175906
transform 1 0 9744 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1538_
timestamp 1698175906
transform -1 0 10416 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1539_
timestamp 1698175906
transform 1 0 5936 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1540_
timestamp 1698175906
transform -1 0 6720 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698175906
transform 1 0 7616 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1542_
timestamp 1698175906
transform 1 0 6720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1698175906
transform -1 0 5488 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1544_
timestamp 1698175906
transform -1 0 5600 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1545_
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1546_
timestamp 1698175906
transform 1 0 5488 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1547_
timestamp 1698175906
transform -1 0 7168 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1548_
timestamp 1698175906
transform -1 0 7728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1549_
timestamp 1698175906
transform 1 0 6496 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1550_
timestamp 1698175906
transform -1 0 7280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1551_
timestamp 1698175906
transform 1 0 19824 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1552_
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1553_
timestamp 1698175906
transform 1 0 9184 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1554_
timestamp 1698175906
transform 1 0 5264 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1555_
timestamp 1698175906
transform 1 0 5600 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1556_
timestamp 1698175906
transform -1 0 7168 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1557_
timestamp 1698175906
transform 1 0 6384 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1558_
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1559_
timestamp 1698175906
transform -1 0 3136 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1560_
timestamp 1698175906
transform 1 0 4816 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1698175906
transform 1 0 5712 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1698175906
transform 1 0 6384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1563_
timestamp 1698175906
transform -1 0 7952 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1564_
timestamp 1698175906
transform -1 0 11536 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1565_
timestamp 1698175906
transform -1 0 7168 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1566_
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1567_
timestamp 1698175906
transform 1 0 6384 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1568_
timestamp 1698175906
transform -1 0 6384 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1569_
timestamp 1698175906
transform 1 0 6496 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1570_
timestamp 1698175906
transform -1 0 6496 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1571_
timestamp 1698175906
transform 1 0 6048 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1572_
timestamp 1698175906
transform 1 0 4592 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1573_
timestamp 1698175906
transform 1 0 5488 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1574_
timestamp 1698175906
transform -1 0 7056 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1575_
timestamp 1698175906
transform 1 0 5600 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1576_
timestamp 1698175906
transform 1 0 5376 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1577_
timestamp 1698175906
transform 1 0 6384 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1578_
timestamp 1698175906
transform 1 0 8064 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1579_
timestamp 1698175906
transform 1 0 8736 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1580_
timestamp 1698175906
transform -1 0 7616 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1581_
timestamp 1698175906
transform -1 0 6048 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1582_
timestamp 1698175906
transform -1 0 6944 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1583_
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1584_
timestamp 1698175906
transform -1 0 3248 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1585_
timestamp 1698175906
transform 1 0 4704 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1586_
timestamp 1698175906
transform -1 0 6496 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1587_
timestamp 1698175906
transform -1 0 3136 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1588_
timestamp 1698175906
transform -1 0 9856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1698175906
transform 1 0 7280 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1590_
timestamp 1698175906
transform -1 0 9744 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1591_
timestamp 1698175906
transform 1 0 7840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1592_
timestamp 1698175906
transform -1 0 10864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1593_
timestamp 1698175906
transform 1 0 9856 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1594_
timestamp 1698175906
transform 1 0 12544 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1595_
timestamp 1698175906
transform 1 0 10864 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1596_
timestamp 1698175906
transform -1 0 14560 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1698175906
transform -1 0 40208 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1698175906
transform -1 0 39984 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1698175906
transform -1 0 45920 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1600_
timestamp 1698175906
transform -1 0 45472 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1601_
timestamp 1698175906
transform -1 0 45584 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1602_
timestamp 1698175906
transform 1 0 3360 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1603_
timestamp 1698175906
transform 1 0 30800 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1604_
timestamp 1698175906
transform -1 0 26432 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1605_
timestamp 1698175906
transform -1 0 26880 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1606_
timestamp 1698175906
transform 1 0 24640 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1607_
timestamp 1698175906
transform -1 0 20944 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1698175906
transform -1 0 20048 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1609_
timestamp 1698175906
transform -1 0 24416 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1610_
timestamp 1698175906
transform -1 0 23744 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1611_
timestamp 1698175906
transform -1 0 20832 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1612_
timestamp 1698175906
transform -1 0 23744 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1613_
timestamp 1698175906
transform -1 0 18928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1614_
timestamp 1698175906
transform -1 0 27216 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1615_
timestamp 1698175906
transform -1 0 22960 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1616_
timestamp 1698175906
transform -1 0 19712 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1617_
timestamp 1698175906
transform -1 0 23184 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1618_
timestamp 1698175906
transform -1 0 21840 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1619_
timestamp 1698175906
transform -1 0 24864 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1620_
timestamp 1698175906
transform 1 0 24864 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1621_
timestamp 1698175906
transform 1 0 27104 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1622_
timestamp 1698175906
transform 1 0 28000 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698175906
transform -1 0 10192 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1624_
timestamp 1698175906
transform 1 0 8736 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1626_
timestamp 1698175906
transform 1 0 35728 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698175906
transform -1 0 38304 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1628_
timestamp 1698175906
transform 1 0 30240 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1629_
timestamp 1698175906
transform -1 0 37744 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1630_
timestamp 1698175906
transform -1 0 34720 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698175906
transform 1 0 33376 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1632_
timestamp 1698175906
transform 1 0 33712 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1698175906
transform -1 0 35280 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698175906
transform 1 0 33264 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1635_
timestamp 1698175906
transform 1 0 33600 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1636_
timestamp 1698175906
transform 1 0 40208 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698175906
transform 1 0 40992 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1638_
timestamp 1698175906
transform 1 0 40768 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1639_
timestamp 1698175906
transform -1 0 42224 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1640_
timestamp 1698175906
transform -1 0 41776 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1641_
timestamp 1698175906
transform -1 0 45808 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1642_
timestamp 1698175906
transform 1 0 43904 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1643_
timestamp 1698175906
transform 1 0 37632 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1644_
timestamp 1698175906
transform 1 0 44688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1645_
timestamp 1698175906
transform 1 0 45808 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1698175906
transform 1 0 44688 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1647_
timestamp 1698175906
transform 1 0 44912 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1648_
timestamp 1698175906
transform -1 0 45248 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1698175906
transform 1 0 44800 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1650_
timestamp 1698175906
transform -1 0 44800 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1651_
timestamp 1698175906
transform 1 0 39648 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1698175906
transform 1 0 39984 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1653_
timestamp 1698175906
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1654_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44688 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1655_
timestamp 1698175906
transform 1 0 45696 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1656_
timestamp 1698175906
transform 1 0 47936 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1657_
timestamp 1698175906
transform 1 0 50176 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1658_
timestamp 1698175906
transform 1 0 50176 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1659_
timestamp 1698175906
transform -1 0 53424 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1660_
timestamp 1698175906
transform -1 0 53424 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1661_
timestamp 1698175906
transform 1 0 45136 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1662_
timestamp 1698175906
transform 1 0 50176 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1663_
timestamp 1698175906
transform 1 0 50176 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1664_
timestamp 1698175906
transform 1 0 46480 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1665_
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1666_
timestamp 1698175906
transform 1 0 46032 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1667_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1668_
timestamp 1698175906
transform 1 0 30688 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1669_
timestamp 1698175906
transform 1 0 30576 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1670_
timestamp 1698175906
transform 1 0 29456 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1671_
timestamp 1698175906
transform -1 0 44464 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1672_
timestamp 1698175906
transform -1 0 44912 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1673_
timestamp 1698175906
transform 1 0 33824 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1674_
timestamp 1698175906
transform 1 0 35280 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1675_
timestamp 1698175906
transform 1 0 37856 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1676_
timestamp 1698175906
transform 1 0 40992 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1677_
timestamp 1698175906
transform 1 0 26656 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1678_
timestamp 1698175906
transform 1 0 26432 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1679_
timestamp 1698175906
transform -1 0 24864 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1680_
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1681_
timestamp 1698175906
transform 1 0 20720 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1682_
timestamp 1698175906
transform 1 0 20384 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1683_
timestamp 1698175906
transform 1 0 20496 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1684_
timestamp 1698175906
transform 1 0 24080 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1685_
timestamp 1698175906
transform 1 0 31024 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1686_
timestamp 1698175906
transform 1 0 31024 0 1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1687_
timestamp 1698175906
transform -1 0 30016 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1688_
timestamp 1698175906
transform -1 0 32592 0 1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1689_
timestamp 1698175906
transform 1 0 31248 0 1 28224
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1690_
timestamp 1698175906
transform 1 0 33824 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1691_
timestamp 1698175906
transform 1 0 32816 0 1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1692_
timestamp 1698175906
transform 1 0 35168 0 -1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1693_
timestamp 1698175906
transform 1 0 35168 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1694_
timestamp 1698175906
transform 1 0 50176 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1695_
timestamp 1698175906
transform -1 0 53424 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1696_
timestamp 1698175906
transform 1 0 45808 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1697_
timestamp 1698175906
transform 1 0 46368 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1698_
timestamp 1698175906
transform -1 0 53424 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1699_
timestamp 1698175906
transform 1 0 50176 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1700_
timestamp 1698175906
transform 1 0 50176 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1701_
timestamp 1698175906
transform 1 0 50176 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1702_
timestamp 1698175906
transform 1 0 50176 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1703_
timestamp 1698175906
transform 1 0 45584 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1704_
timestamp 1698175906
transform 1 0 50176 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1705_
timestamp 1698175906
transform 1 0 50176 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1706_
timestamp 1698175906
transform 1 0 46928 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1707_
timestamp 1698175906
transform -1 0 52192 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1708_
timestamp 1698175906
transform -1 0 25760 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1709_
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1710_
timestamp 1698175906
transform 1 0 26880 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1711_
timestamp 1698175906
transform -1 0 28000 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1712_
timestamp 1698175906
transform -1 0 21392 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1713_
timestamp 1698175906
transform 1 0 20720 0 -1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1714_
timestamp 1698175906
transform -1 0 23296 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1715_
timestamp 1698175906
transform 1 0 22960 0 1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1716_
timestamp 1698175906
transform 1 0 31696 0 1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1717_
timestamp 1698175906
transform 1 0 35280 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1718_
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1719_
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1720_
timestamp 1698175906
transform 1 0 39648 0 1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1721_
timestamp 1698175906
transform 1 0 35728 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1722_
timestamp 1698175906
transform -1 0 44016 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1723_
timestamp 1698175906
transform 1 0 41776 0 -1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1724_
timestamp 1698175906
transform 1 0 26096 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1725_
timestamp 1698175906
transform 1 0 18032 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1726_
timestamp 1698175906
transform 1 0 21840 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1727_
timestamp 1698175906
transform 1 0 15232 0 1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1728_
timestamp 1698175906
transform 1 0 16688 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1729_
timestamp 1698175906
transform -1 0 31024 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1730_
timestamp 1698175906
transform -1 0 32256 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1731_
timestamp 1698175906
transform -1 0 32368 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1732_
timestamp 1698175906
transform 1 0 25424 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1733_
timestamp 1698175906
transform 1 0 16016 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1734_
timestamp 1698175906
transform 1 0 14560 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1735_
timestamp 1698175906
transform 1 0 12768 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1736_
timestamp 1698175906
transform 1 0 6608 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1737_
timestamp 1698175906
transform 1 0 9520 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1738_
timestamp 1698175906
transform 1 0 7168 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1739_
timestamp 1698175906
transform 1 0 11872 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1740_
timestamp 1698175906
transform 1 0 31696 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1741_
timestamp 1698175906
transform 1 0 32256 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1742_
timestamp 1698175906
transform -1 0 40096 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1743_
timestamp 1698175906
transform -1 0 43344 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1744_
timestamp 1698175906
transform 1 0 42560 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1745_
timestamp 1698175906
transform 1 0 43232 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1746_
timestamp 1698175906
transform 1 0 41216 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1747_
timestamp 1698175906
transform 1 0 37296 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1748_
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1749_
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1750_
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1751_
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1752_
timestamp 1698175906
transform -1 0 5264 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1753_
timestamp 1698175906
transform 1 0 5152 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1754_
timestamp 1698175906
transform 1 0 7168 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1755_
timestamp 1698175906
transform 1 0 10080 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1756_
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1757_
timestamp 1698175906
transform 1 0 14448 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1758_
timestamp 1698175906
transform 1 0 16464 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1759_
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1760_
timestamp 1698175906
transform 1 0 17696 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1761_
timestamp 1698175906
transform 1 0 12320 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1762_
timestamp 1698175906
transform 1 0 9408 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1763_
timestamp 1698175906
transform 1 0 13216 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1764_
timestamp 1698175906
transform 1 0 9632 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1765_
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1766_
timestamp 1698175906
transform 1 0 13776 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1767_
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1768_
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1769_
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1770_
timestamp 1698175906
transform 1 0 5488 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1771_
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1772_
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1773_
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1774_
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1775_
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1776_
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1777_
timestamp 1698175906
transform 1 0 9856 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1778_
timestamp 1698175906
transform 1 0 13328 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1779_
timestamp 1698175906
transform 1 0 45472 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1780_
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1781_
timestamp 1698175906
transform -1 0 29680 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1782_
timestamp 1698175906
transform 1 0 19824 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1783_
timestamp 1698175906
transform 1 0 19488 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1784_
timestamp 1698175906
transform 1 0 16800 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1785_
timestamp 1698175906
transform 1 0 15792 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1786_
timestamp 1698175906
transform 1 0 19824 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1787_
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1788_
timestamp 1698175906
transform -1 0 30912 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1789_
timestamp 1698175906
transform 1 0 8848 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1790_
timestamp 1698175906
transform 1 0 35728 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1791_
timestamp 1698175906
transform 1 0 29456 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1792_
timestamp 1698175906
transform 1 0 30128 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1793_
timestamp 1698175906
transform 1 0 39984 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1794_
timestamp 1698175906
transform -1 0 47712 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1795_
timestamp 1698175906
transform -1 0 49504 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1796_
timestamp 1698175906
transform 1 0 42784 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1797_
timestamp 1698175906
transform -1 0 42336 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__I
timestamp 1698175906
transform -1 0 39872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__I
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__A1
timestamp 1698175906
transform 1 0 44912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__B2
timestamp 1698175906
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__A1
timestamp 1698175906
transform -1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A1
timestamp 1698175906
transform 1 0 40992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__B2
timestamp 1698175906
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A1
timestamp 1698175906
transform -1 0 35392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__I
timestamp 1698175906
transform 1 0 44912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__I
timestamp 1698175906
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__A2
timestamp 1698175906
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1698175906
transform 1 0 44912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A2
timestamp 1698175906
transform 1 0 45360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698175906
transform 1 0 39200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__I
timestamp 1698175906
transform 1 0 38080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1698175906
transform 1 0 47376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I
timestamp 1698175906
transform -1 0 45584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A1
timestamp 1698175906
transform 1 0 46032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698175906
transform 1 0 45920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__I
timestamp 1698175906
transform -1 0 31024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__I
timestamp 1698175906
transform 1 0 48048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698175906
transform -1 0 47152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A2
timestamp 1698175906
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A2
timestamp 1698175906
transform 1 0 51184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__A2
timestamp 1698175906
transform 1 0 51744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698175906
transform 1 0 51296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0901__A2
timestamp 1698175906
transform 1 0 49840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698175906
transform 1 0 52080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A2
timestamp 1698175906
transform 1 0 50176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A1
timestamp 1698175906
transform 1 0 51184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A1
timestamp 1698175906
transform 1 0 48160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A2
timestamp 1698175906
transform 1 0 49392 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A1
timestamp 1698175906
transform 1 0 46256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A3
timestamp 1698175906
transform 1 0 43232 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__I
timestamp 1698175906
transform 1 0 44912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A2
timestamp 1698175906
transform 1 0 42784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__A1
timestamp 1698175906
transform 1 0 46032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__I
timestamp 1698175906
transform -1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1698175906
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A1
timestamp 1698175906
transform 1 0 29792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A2
timestamp 1698175906
transform 1 0 30240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A1
timestamp 1698175906
transform 1 0 26544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__A1
timestamp 1698175906
transform -1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__A2
timestamp 1698175906
transform 1 0 42784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__C
timestamp 1698175906
transform 1 0 31024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__A2
timestamp 1698175906
transform 1 0 37520 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__I
timestamp 1698175906
transform 1 0 44912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__B
timestamp 1698175906
transform 1 0 30912 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__I
timestamp 1698175906
transform 1 0 26096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__C
timestamp 1698175906
transform 1 0 31136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A1
timestamp 1698175906
transform 1 0 42672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A1
timestamp 1698175906
transform 1 0 43008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__B
timestamp 1698175906
transform 1 0 36288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__B
timestamp 1698175906
transform -1 0 36176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__B
timestamp 1698175906
transform -1 0 37968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__B
timestamp 1698175906
transform -1 0 43120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A2
timestamp 1698175906
transform 1 0 43792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A3
timestamp 1698175906
transform -1 0 43792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__C
timestamp 1698175906
transform -1 0 28000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I
timestamp 1698175906
transform 1 0 29344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__B
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1015__B
timestamp 1698175906
transform 1 0 24304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__I
timestamp 1698175906
transform 1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__I
timestamp 1698175906
transform 1 0 30688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__I
timestamp 1698175906
transform 1 0 26096 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__B
timestamp 1698175906
transform -1 0 27664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A1
timestamp 1698175906
transform -1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__I0
timestamp 1698175906
transform 1 0 34160 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698175906
transform 1 0 43344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A2
timestamp 1698175906
transform -1 0 44912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__I
timestamp 1698175906
transform 1 0 30352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__I
timestamp 1698175906
transform 1 0 45024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A1
timestamp 1698175906
transform 1 0 32704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__I
timestamp 1698175906
transform 1 0 34496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I
timestamp 1698175906
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698175906
transform 1 0 32144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698175906
transform 1 0 30464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698175906
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__I
timestamp 1698175906
transform 1 0 35504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698175906
transform 1 0 31808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A1
timestamp 1698175906
transform 1 0 32256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698175906
transform -1 0 32032 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A1
timestamp 1698175906
transform 1 0 32144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__I
timestamp 1698175906
transform 1 0 35728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698175906
transform 1 0 35280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__A1
timestamp 1698175906
transform 1 0 33824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698175906
transform 1 0 34832 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698175906
transform -1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698175906
transform 1 0 35952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698175906
transform -1 0 35504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698175906
transform 1 0 35504 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A1
timestamp 1698175906
transform 1 0 34608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A2
timestamp 1698175906
transform 1 0 47600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A3
timestamp 1698175906
transform 1 0 48944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__I
timestamp 1698175906
transform -1 0 49504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698175906
transform 1 0 43232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__I
timestamp 1698175906
transform 1 0 43904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698175906
transform 1 0 38304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__A2
timestamp 1698175906
transform 1 0 45360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__I
timestamp 1698175906
transform 1 0 28784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__B1
timestamp 1698175906
transform 1 0 42112 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__B2
timestamp 1698175906
transform 1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__I
timestamp 1698175906
transform 1 0 42784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698175906
transform 1 0 30352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698175906
transform 1 0 43792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A2
timestamp 1698175906
transform 1 0 42560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__B2
timestamp 1698175906
transform -1 0 34384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A2
timestamp 1698175906
transform 1 0 45584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A1
timestamp 1698175906
transform 1 0 49840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698175906
transform 1 0 29456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__B1
timestamp 1698175906
transform 1 0 29008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__B2
timestamp 1698175906
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A1
timestamp 1698175906
transform 1 0 37744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__B2
timestamp 1698175906
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__I
timestamp 1698175906
transform 1 0 44240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__B
timestamp 1698175906
transform 1 0 48832 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A2
timestamp 1698175906
transform -1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A1
timestamp 1698175906
transform 1 0 30128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__B1
timestamp 1698175906
transform 1 0 29680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__B2
timestamp 1698175906
transform 1 0 30576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A1
timestamp 1698175906
transform -1 0 37968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__B2
timestamp 1698175906
transform -1 0 43680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__B
timestamp 1698175906
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A2
timestamp 1698175906
transform 1 0 45248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__I
timestamp 1698175906
transform -1 0 30352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__B1
timestamp 1698175906
transform 1 0 29232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A1
timestamp 1698175906
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__B2
timestamp 1698175906
transform -1 0 37296 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698175906
transform 1 0 51632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__I
timestamp 1698175906
transform 1 0 28000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A1
timestamp 1698175906
transform -1 0 38752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__B2
timestamp 1698175906
transform -1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A3
timestamp 1698175906
transform -1 0 41776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698175906
transform -1 0 50736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__I
timestamp 1698175906
transform 1 0 30688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__I
timestamp 1698175906
transform 1 0 48496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__A1
timestamp 1698175906
transform 1 0 37856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A3
timestamp 1698175906
transform 1 0 42560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A1
timestamp 1698175906
transform -1 0 39648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__B2
timestamp 1698175906
transform -1 0 41104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698175906
transform 1 0 44800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A3
timestamp 1698175906
transform 1 0 43344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__B2
timestamp 1698175906
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__A1
timestamp 1698175906
transform 1 0 38416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__B2
timestamp 1698175906
transform -1 0 39872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A1
timestamp 1698175906
transform -1 0 43008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A3
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A2
timestamp 1698175906
transform -1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A2
timestamp 1698175906
transform -1 0 19712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A2
timestamp 1698175906
transform -1 0 21504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A2
timestamp 1698175906
transform 1 0 15680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A2
timestamp 1698175906
transform -1 0 29904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A2
timestamp 1698175906
transform 1 0 27216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__A2
timestamp 1698175906
transform 1 0 29232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A2
timestamp 1698175906
transform -1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__A1
timestamp 1698175906
transform -1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__A2
timestamp 1698175906
transform 1 0 27104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A2
timestamp 1698175906
transform -1 0 23520 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A2
timestamp 1698175906
transform 1 0 24192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__A2
timestamp 1698175906
transform -1 0 23072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1181__A2
timestamp 1698175906
transform -1 0 31696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A2
timestamp 1698175906
transform 1 0 46816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__I
timestamp 1698175906
transform -1 0 39536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1186__A2
timestamp 1698175906
transform -1 0 46032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__B
timestamp 1698175906
transform 1 0 45920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__A3
timestamp 1698175906
transform 1 0 48160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__B
timestamp 1698175906
transform -1 0 49280 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1198__A1
timestamp 1698175906
transform 1 0 47488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__A1
timestamp 1698175906
transform -1 0 46928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__A1
timestamp 1698175906
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__I0
timestamp 1698175906
transform 1 0 48048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698175906
transform 1 0 46480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A1
timestamp 1698175906
transform -1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A2
timestamp 1698175906
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A1
timestamp 1698175906
transform 1 0 25536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A1
timestamp 1698175906
transform 1 0 27104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__C
timestamp 1698175906
transform -1 0 27552 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__A1
timestamp 1698175906
transform 1 0 30688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__A1
timestamp 1698175906
transform 1 0 30240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__C
timestamp 1698175906
transform -1 0 28224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1213__A1
timestamp 1698175906
transform 1 0 28112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__A2
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698175906
transform 1 0 25984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__B
timestamp 1698175906
transform 1 0 26656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1218__A1
timestamp 1698175906
transform -1 0 27104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__B
timestamp 1698175906
transform 1 0 26992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A1
timestamp 1698175906
transform 1 0 23072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698175906
transform 1 0 21504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1229__A1
timestamp 1698175906
transform 1 0 22736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__A1
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__A1
timestamp 1698175906
transform 1 0 23184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__A1
timestamp 1698175906
transform 1 0 35168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__A1
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__A1
timestamp 1698175906
transform 1 0 34272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698175906
transform 1 0 33152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A1
timestamp 1698175906
transform 1 0 41328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1249__A1
timestamp 1698175906
transform 1 0 41776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__B
timestamp 1698175906
transform 1 0 40544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A1
timestamp 1698175906
transform 1 0 35840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__B
timestamp 1698175906
transform -1 0 36848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698175906
transform 1 0 40992 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__B
timestamp 1698175906
transform 1 0 41440 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__A1
timestamp 1698175906
transform 1 0 40992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698175906
transform 1 0 38976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__B
timestamp 1698175906
transform 1 0 39424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__I
timestamp 1698175906
transform 1 0 31696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__I
timestamp 1698175906
transform 1 0 28784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__I
timestamp 1698175906
transform 1 0 32704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698175906
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__A2
timestamp 1698175906
transform 1 0 25984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__A2
timestamp 1698175906
transform -1 0 26208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__B
timestamp 1698175906
transform -1 0 26432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__I
timestamp 1698175906
transform 1 0 15120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A1
timestamp 1698175906
transform 1 0 21952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__C
timestamp 1698175906
transform 1 0 19600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698175906
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__B
timestamp 1698175906
transform -1 0 24640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__I
timestamp 1698175906
transform -1 0 18592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__B
timestamp 1698175906
transform -1 0 27216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__A1
timestamp 1698175906
transform 1 0 28000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__I
timestamp 1698175906
transform 1 0 26320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698175906
transform 1 0 26320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__B
timestamp 1698175906
transform 1 0 24080 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__B
timestamp 1698175906
transform 1 0 16800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698175906
transform -1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698175906
transform -1 0 16016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__B
timestamp 1698175906
transform 1 0 14784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__I
timestamp 1698175906
transform 1 0 11648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__I
timestamp 1698175906
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__B
timestamp 1698175906
transform 1 0 10416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__B
timestamp 1698175906
transform 1 0 11424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A2
timestamp 1698175906
transform 1 0 11648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__B
timestamp 1698175906
transform 1 0 10864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__B
timestamp 1698175906
transform -1 0 14896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__I
timestamp 1698175906
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__C
timestamp 1698175906
transform -1 0 14672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A1
timestamp 1698175906
transform 1 0 38304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__I
timestamp 1698175906
transform -1 0 42336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__I
timestamp 1698175906
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A1
timestamp 1698175906
transform 1 0 41216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A1
timestamp 1698175906
transform 1 0 41888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__B
timestamp 1698175906
transform 1 0 36176 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A2
timestamp 1698175906
transform 1 0 31472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A1
timestamp 1698175906
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698175906
transform 1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698175906
transform 1 0 17248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__A2
timestamp 1698175906
transform -1 0 17024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__A2
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A1
timestamp 1698175906
transform 1 0 13104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A2
timestamp 1698175906
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A2
timestamp 1698175906
transform 1 0 14000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A2
timestamp 1698175906
transform 1 0 12432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__I
timestamp 1698175906
transform 1 0 9072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A2
timestamp 1698175906
transform 1 0 20160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A2
timestamp 1698175906
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A2
timestamp 1698175906
transform 1 0 18704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698175906
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1698175906
transform -1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__A2
timestamp 1698175906
transform 1 0 19040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A2
timestamp 1698175906
transform 1 0 18816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A1
timestamp 1698175906
transform -1 0 32928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698175906
transform 1 0 9632 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1427__A1
timestamp 1698175906
transform -1 0 11200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A1
timestamp 1698175906
transform 1 0 9632 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1698175906
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__C
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__I
timestamp 1698175906
transform -1 0 10864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__B
timestamp 1698175906
transform 1 0 7504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__A1
timestamp 1698175906
transform 1 0 10640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__C
timestamp 1698175906
transform 1 0 7392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__B
timestamp 1698175906
transform -1 0 10528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A1
timestamp 1698175906
transform -1 0 12320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A2
timestamp 1698175906
transform 1 0 13104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__C
timestamp 1698175906
transform -1 0 12208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A1
timestamp 1698175906
transform -1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__C
timestamp 1698175906
transform -1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__A1
timestamp 1698175906
transform 1 0 14560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__C
timestamp 1698175906
transform 1 0 15344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__A1
timestamp 1698175906
transform 1 0 16800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A1
timestamp 1698175906
transform 1 0 19040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A1
timestamp 1698175906
transform 1 0 19040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__A1
timestamp 1698175906
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__A1
timestamp 1698175906
transform -1 0 15904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A1
timestamp 1698175906
transform -1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__I
timestamp 1698175906
transform 1 0 10528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A1
timestamp 1698175906
transform 1 0 13328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1698175906
transform 1 0 8624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A1
timestamp 1698175906
transform 1 0 10640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A1
timestamp 1698175906
transform -1 0 3584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__I
timestamp 1698175906
transform 1 0 11536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__B
timestamp 1698175906
transform -1 0 8400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__B
timestamp 1698175906
transform 1 0 7168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__B
timestamp 1698175906
transform 1 0 7504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__I
timestamp 1698175906
transform 1 0 5152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A1
timestamp 1698175906
transform 1 0 3472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A1
timestamp 1698175906
transform -1 0 4704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A1
timestamp 1698175906
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A1
timestamp 1698175906
transform 1 0 3360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A1
timestamp 1698175906
transform 1 0 7056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__C
timestamp 1698175906
transform 1 0 14784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A1
timestamp 1698175906
transform 1 0 45920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A1
timestamp 1698175906
transform 1 0 45696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A1
timestamp 1698175906
transform -1 0 44464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__B
timestamp 1698175906
transform 1 0 43792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698175906
transform -1 0 31920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1698175906
transform 1 0 25424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__C
timestamp 1698175906
transform -1 0 27328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A1
timestamp 1698175906
transform 1 0 21392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A1
timestamp 1698175906
transform 1 0 25760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A1
timestamp 1698175906
transform 1 0 27776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A1
timestamp 1698175906
transform -1 0 10640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1698175906
transform -1 0 10416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1698175906
transform 1 0 38528 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__I
timestamp 1698175906
transform 1 0 30016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A2
timestamp 1698175906
transform 1 0 34160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1698175906
transform -1 0 34496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1698175906
transform 1 0 37408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__CLK
timestamp 1698175906
transform 1 0 47936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__CLK
timestamp 1698175906
transform 1 0 49168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__CLK
timestamp 1698175906
transform 1 0 51408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__CLK
timestamp 1698175906
transform 1 0 49168 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__CLK
timestamp 1698175906
transform -1 0 50512 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__CLK
timestamp 1698175906
transform 1 0 50848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__CLK
timestamp 1698175906
transform 1 0 49952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__CLK
timestamp 1698175906
transform 1 0 48384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__CLK
timestamp 1698175906
transform 1 0 49952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__CLK
timestamp 1698175906
transform 1 0 49952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__CLK
timestamp 1698175906
transform 1 0 49952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__CLK
timestamp 1698175906
transform -1 0 42112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__CLK
timestamp 1698175906
transform 1 0 49504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__CLK
timestamp 1698175906
transform 1 0 28448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__CLK
timestamp 1698175906
transform 1 0 44688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__CLK
timestamp 1698175906
transform 1 0 45136 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__CLK
timestamp 1698175906
transform 1 0 37296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__CLK
timestamp 1698175906
transform 1 0 38752 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__CLK
timestamp 1698175906
transform 1 0 41328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__CLK
timestamp 1698175906
transform 1 0 44464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__CLK
timestamp 1698175906
transform 1 0 24864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__CLK
timestamp 1698175906
transform 1 0 23968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__CLK
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__CLK
timestamp 1698175906
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__CLK
timestamp 1698175906
transform 1 0 27328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__CLK
timestamp 1698175906
transform 1 0 34720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__CLK
timestamp 1698175906
transform 1 0 30240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__CLK
timestamp 1698175906
transform 1 0 32816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__CLK
timestamp 1698175906
transform 1 0 34944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__CLK
timestamp 1698175906
transform -1 0 37744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__CLK
timestamp 1698175906
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__CLK
timestamp 1698175906
transform 1 0 38864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__CLK
timestamp 1698175906
transform 1 0 38864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__CLK
timestamp 1698175906
transform 1 0 48832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__CLK
timestamp 1698175906
transform 1 0 49952 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__CLK
timestamp 1698175906
transform -1 0 49280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__CLK
timestamp 1698175906
transform 1 0 46144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__CLK
timestamp 1698175906
transform 1 0 50176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__CLK
timestamp 1698175906
transform 1 0 49952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__CLK
timestamp 1698175906
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__CLK
timestamp 1698175906
transform 1 0 49952 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__CLK
timestamp 1698175906
transform 1 0 49952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__CLK
timestamp 1698175906
transform 1 0 46704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__CLK
timestamp 1698175906
transform 1 0 52416 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__CLK
timestamp 1698175906
transform 1 0 25984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__CLK
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__CLK
timestamp 1698175906
transform 1 0 30576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__CLK
timestamp 1698175906
transform 1 0 28224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__CLK
timestamp 1698175906
transform 1 0 17696 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__CLK
timestamp 1698175906
transform 1 0 20496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__CLK
timestamp 1698175906
transform -1 0 23744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__CLK
timestamp 1698175906
transform 1 0 22736 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__CLK
timestamp 1698175906
transform 1 0 31472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__CLK
timestamp 1698175906
transform 1 0 38752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__CLK
timestamp 1698175906
transform -1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__CLK
timestamp 1698175906
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__CLK
timestamp 1698175906
transform 1 0 43344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__CLK
timestamp 1698175906
transform 1 0 39200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__CLK
timestamp 1698175906
transform 1 0 44240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__CLK
timestamp 1698175906
transform 1 0 45472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__CLK
timestamp 1698175906
transform 1 0 29792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__CLK
timestamp 1698175906
transform 1 0 17808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__CLK
timestamp 1698175906
transform 1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__CLK
timestamp 1698175906
transform 1 0 18928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__CLK
timestamp 1698175906
transform 1 0 20160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__CLK
timestamp 1698175906
transform 1 0 31248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__CLK
timestamp 1698175906
transform -1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__CLK
timestamp 1698175906
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__CLK
timestamp 1698175906
transform 1 0 29568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__CLK
timestamp 1698175906
transform 1 0 19264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__CLK
timestamp 1698175906
transform 1 0 18032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__CLK
timestamp 1698175906
transform 1 0 17920 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__CLK
timestamp 1698175906
transform 1 0 10080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__CLK
timestamp 1698175906
transform 1 0 9296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__CLK
timestamp 1698175906
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__CLK
timestamp 1698175906
transform 1 0 35168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__CLK
timestamp 1698175906
transform 1 0 35728 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__CLK
timestamp 1698175906
transform 1 0 44464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__CLK
timestamp 1698175906
transform 1 0 37968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__CLK
timestamp 1698175906
transform -1 0 32480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__CLK
timestamp 1698175906
transform 1 0 4816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__CLK
timestamp 1698175906
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__CLK
timestamp 1698175906
transform 1 0 5712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__CLK
timestamp 1698175906
transform 1 0 8400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__CLK
timestamp 1698175906
transform 1 0 10640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__CLK
timestamp 1698175906
transform 1 0 13552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__CLK
timestamp 1698175906
transform 1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__CLK
timestamp 1698175906
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__CLK
timestamp 1698175906
transform 1 0 22064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__CLK
timestamp 1698175906
transform 1 0 17472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__CLK
timestamp 1698175906
transform 1 0 16240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__CLK
timestamp 1698175906
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__CLK
timestamp 1698175906
transform 1 0 16464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__CLK
timestamp 1698175906
transform 1 0 9408 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__CLK
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__CLK
timestamp 1698175906
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__CLK
timestamp 1698175906
transform -1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__CLK
timestamp 1698175906
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__CLK
timestamp 1698175906
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__CLK
timestamp 1698175906
transform 1 0 8960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__CLK
timestamp 1698175906
transform 1 0 4816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__CLK
timestamp 1698175906
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__CLK
timestamp 1698175906
transform -1 0 5264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__CLK
timestamp 1698175906
transform -1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__CLK
timestamp 1698175906
transform 1 0 4816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__CLK
timestamp 1698175906
transform 1 0 9632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__CLK
timestamp 1698175906
transform 1 0 48944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__CLK
timestamp 1698175906
transform -1 0 16352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__D
timestamp 1698175906
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__CLK
timestamp 1698175906
transform 1 0 19600 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__CLK
timestamp 1698175906
transform 1 0 19264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__CLK
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__CLK
timestamp 1698175906
transform 1 0 15568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__CLK
timestamp 1698175906
transform 1 0 19600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__CLK
timestamp 1698175906
transform 1 0 12320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__CLK
timestamp 1698175906
transform 1 0 39200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__CLK
timestamp 1698175906
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__CLK
timestamp 1698175906
transform 1 0 33376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__CLK
timestamp 1698175906
transform 1 0 43456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__CLK
timestamp 1698175906
transform 1 0 47936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__CLK
timestamp 1698175906
transform 1 0 46032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__CLK
timestamp 1698175906
transform 1 0 46256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__CLK
timestamp 1698175906
transform 1 0 42560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 17696 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 28224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 27104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 9632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 10976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 17920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 18144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 37968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 38528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 47824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 47712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 34832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 34720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 43680 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 52528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 53424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 53424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 52752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 52752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform 1 0 53200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform -1 0 53424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 53424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform -1 0 2800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform -1 0 41328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1698175906
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1698175906
transform -1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1698175906
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27104 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698175906
transform 1 0 14560 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698175906
transform -1 0 26320 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698175906
transform -1 0 8960 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698175906
transform 1 0 6832 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698175906
transform -1 0 17696 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698175906
transform 1 0 15008 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698175906
transform -1 0 43904 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698175906
transform 1 0 39424 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698175906
transform 1 0 48048 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698175906
transform 1 0 47936 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698175906
transform -1 0 37968 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698175906
transform 1 0 34720 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698175906
transform -1 0 47600 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698175906
transform -1 0 46816 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_19
timestamp 1698175906
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_27 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_31 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698175906
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_96
timestamp 1698175906
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_100
timestamp 1698175906
transform 1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_142 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_158
timestamp 1698175906
transform 1 0 19040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_166
timestamp 1698175906
transform 1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_177
timestamp 1698175906
transform 1 0 21168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_193
timestamp 1698175906
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698175906
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698175906
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_235
timestamp 1698175906
transform 1 0 27664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698175906
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_248
timestamp 1698175906
transform 1 0 29120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_252
timestamp 1698175906
transform 1 0 29568 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_257
timestamp 1698175906
transform 1 0 30128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_265
timestamp 1698175906
transform 1 0 31024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698175906
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290
timestamp 1698175906
transform 1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_298
timestamp 1698175906
transform 1 0 34720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_302
timestamp 1698175906
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_334
timestamp 1698175906
transform 1 0 38752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_350
timestamp 1698175906
transform 1 0 40544 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_358
timestamp 1698175906
transform 1 0 41440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_364
timestamp 1698175906
transform 1 0 42112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698175906
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698175906
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_452
timestamp 1698175906
transform 1 0 51968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_454
timestamp 1698175906
transform 1 0 52192 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_88
timestamp 1698175906
transform 1 0 11200 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_92
timestamp 1698175906
transform 1 0 11648 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_119
timestamp 1698175906
transform 1 0 14672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_123
timestamp 1698175906
transform 1 0 15120 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698175906
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 19040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 19488 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_194
timestamp 1698175906
transform 1 0 23072 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_217
timestamp 1698175906
transform 1 0 25648 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_233
timestamp 1698175906
transform 1 0 27440 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_264
timestamp 1698175906
transform 1 0 30912 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_298
timestamp 1698175906
transform 1 0 34720 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_302
timestamp 1698175906
transform 1 0 35168 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_332
timestamp 1698175906
transform 1 0 38528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_336
timestamp 1698175906
transform 1 0 38976 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_344
timestamp 1698175906
transform 1 0 39872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_383
timestamp 1698175906
transform 1 0 44240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_387
timestamp 1698175906
transform 1 0 44688 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_403
timestamp 1698175906
transform 1 0 46480 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_415
timestamp 1698175906
transform 1 0 47824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698175906
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_426
timestamp 1698175906
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_53
timestamp 1698175906
transform 1 0 7280 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_61
timestamp 1698175906
transform 1 0 8176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_65
timestamp 1698175906
transform 1 0 8624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_96
timestamp 1698175906
transform 1 0 12096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_100
timestamp 1698175906
transform 1 0 12544 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698175906
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_123
timestamp 1698175906
transform 1 0 15120 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_164
timestamp 1698175906
transform 1 0 19712 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_172
timestamp 1698175906
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698175906
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_183
timestamp 1698175906
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_185
timestamp 1698175906
transform 1 0 22064 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_195
timestamp 1698175906
transform 1 0 23184 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_203
timestamp 1698175906
transform 1 0 24080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_207
timestamp 1698175906
transform 1 0 24528 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_209
timestamp 1698175906
transform 1 0 24752 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_216
timestamp 1698175906
transform 1 0 25536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_220
timestamp 1698175906
transform 1 0 25984 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698175906
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_263
timestamp 1698175906
transform 1 0 30800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_294
timestamp 1698175906
transform 1 0 34272 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_310
timestamp 1698175906
transform 1 0 36064 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_314
timestamp 1698175906
transform 1 0 36512 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_325
timestamp 1698175906
transform 1 0 37744 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_355
timestamp 1698175906
transform 1 0 41104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_359
timestamp 1698175906
transform 1 0 41552 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_375
timestamp 1698175906
transform 1 0 43344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_383
timestamp 1698175906
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_391
timestamp 1698175906
transform 1 0 45136 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_399
timestamp 1698175906
transform 1 0 46032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_432
timestamp 1698175906
transform 1 0 49728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_436
timestamp 1698175906
transform 1 0 50176 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698175906
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698175906
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_457
timestamp 1698175906
transform 1 0 52528 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_77
timestamp 1698175906
transform 1 0 9968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_81
timestamp 1698175906
transform 1 0 10416 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_113
timestamp 1698175906
transform 1 0 14000 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_117
timestamp 1698175906
transform 1 0 14448 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_122
timestamp 1698175906
transform 1 0 15008 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_130
timestamp 1698175906
transform 1 0 15904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_134
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_138
timestamp 1698175906
transform 1 0 16800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_174
timestamp 1698175906
transform 1 0 20832 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_182
timestamp 1698175906
transform 1 0 21728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_193
timestamp 1698175906
transform 1 0 22960 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_228
timestamp 1698175906
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_239
timestamp 1698175906
transform 1 0 28112 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_271
timestamp 1698175906
transform 1 0 31696 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698175906
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_319
timestamp 1698175906
transform 1 0 37072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_323
timestamp 1698175906
transform 1 0 37520 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_339
timestamp 1698175906
transform 1 0 39312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698175906
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698175906
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698175906
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_430
timestamp 1698175906
transform 1 0 49504 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_53
timestamp 1698175906
transform 1 0 7280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_61
timestamp 1698175906
transform 1 0 8176 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_65
timestamp 1698175906
transform 1 0 8624 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_79
timestamp 1698175906
transform 1 0 10192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_83
timestamp 1698175906
transform 1 0 10640 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698175906
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698175906
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_136
timestamp 1698175906
transform 1 0 16576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_167
timestamp 1698175906
transform 1 0 20048 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_193
timestamp 1698175906
transform 1 0 22960 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_197
timestamp 1698175906
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_199
timestamp 1698175906
transform 1 0 23632 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_206
timestamp 1698175906
transform 1 0 24416 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_222
timestamp 1698175906
transform 1 0 26208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_224
timestamp 1698175906
transform 1 0 26432 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_231
timestamp 1698175906
transform 1 0 27216 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_239
timestamp 1698175906
transform 1 0 28112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698175906
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_255
timestamp 1698175906
transform 1 0 29904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_257
timestamp 1698175906
transform 1 0 30128 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_270
timestamp 1698175906
transform 1 0 31584 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_274
timestamp 1698175906
transform 1 0 32032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_291
timestamp 1698175906
transform 1 0 33936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_295
timestamp 1698175906
transform 1 0 34384 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_333
timestamp 1698175906
transform 1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_335
timestamp 1698175906
transform 1 0 38864 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_341
timestamp 1698175906
transform 1 0 39536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_349
timestamp 1698175906
transform 1 0 40432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_356
timestamp 1698175906
transform 1 0 41216 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_372
timestamp 1698175906
transform 1 0 43008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_406
timestamp 1698175906
transform 1 0 46816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_427
timestamp 1698175906
transform 1 0 49168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_444
timestamp 1698175906
transform 1 0 51072 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_452
timestamp 1698175906
transform 1 0 51968 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_22
timestamp 1698175906
transform 1 0 3808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_30
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_67
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698175906
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_76
timestamp 1698175906
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_107
timestamp 1698175906
transform 1 0 13328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_111
timestamp 1698175906
transform 1 0 13776 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_127
timestamp 1698175906
transform 1 0 15568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_135
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698175906
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_150
timestamp 1698175906
transform 1 0 18144 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_157
timestamp 1698175906
transform 1 0 18928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_159
timestamp 1698175906
transform 1 0 19152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_200
timestamp 1698175906
transform 1 0 23744 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_208
timestamp 1698175906
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_214
timestamp 1698175906
transform 1 0 25312 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_217
timestamp 1698175906
transform 1 0 25648 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_253
timestamp 1698175906
transform 1 0 29680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_261
timestamp 1698175906
transform 1 0 30576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_269
timestamp 1698175906
transform 1 0 31472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_273
timestamp 1698175906
transform 1 0 31920 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698175906
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698175906
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_298
timestamp 1698175906
transform 1 0 34720 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_306
timestamp 1698175906
transform 1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_308
timestamp 1698175906
transform 1 0 35840 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_319
timestamp 1698175906
transform 1 0 37072 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_323
timestamp 1698175906
transform 1 0 37520 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_369
timestamp 1698175906
transform 1 0 42672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_373
timestamp 1698175906
transform 1 0 43120 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_379
timestamp 1698175906
transform 1 0 43792 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_395
timestamp 1698175906
transform 1 0 45584 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698175906
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_426
timestamp 1698175906
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_440
timestamp 1698175906
transform 1 0 50624 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_448
timestamp 1698175906
transform 1 0 51520 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_452
timestamp 1698175906
transform 1 0 51968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_460
timestamp 1698175906
transform 1 0 52864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_462
timestamp 1698175906
transform 1 0 53088 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_45
timestamp 1698175906
transform 1 0 6384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_49
timestamp 1698175906
transform 1 0 6832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_51
timestamp 1698175906
transform 1 0 7056 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_81
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_85
timestamp 1698175906
transform 1 0 10864 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_115
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_146
timestamp 1698175906
transform 1 0 17696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_150
timestamp 1698175906
transform 1 0 18144 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_158
timestamp 1698175906
transform 1 0 19040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_160
timestamp 1698175906
transform 1 0 19264 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_167
timestamp 1698175906
transform 1 0 20048 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698175906
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_185
timestamp 1698175906
transform 1 0 22064 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_189
timestamp 1698175906
transform 1 0 22512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_200
timestamp 1698175906
transform 1 0 23744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_228
timestamp 1698175906
transform 1 0 26880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_232
timestamp 1698175906
transform 1 0 27328 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_240
timestamp 1698175906
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698175906
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698175906
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698175906
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_261
timestamp 1698175906
transform 1 0 30576 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_291
timestamp 1698175906
transform 1 0 33936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_295
timestamp 1698175906
transform 1 0 34384 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_310
timestamp 1698175906
transform 1 0 36064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698175906
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_323
timestamp 1698175906
transform 1 0 37520 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_331
timestamp 1698175906
transform 1 0 38416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_342
timestamp 1698175906
transform 1 0 39648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_350
timestamp 1698175906
transform 1 0 40544 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_354
timestamp 1698175906
transform 1 0 40992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_356
timestamp 1698175906
transform 1 0 41216 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_363
timestamp 1698175906
transform 1 0 42000 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_367
timestamp 1698175906
transform 1 0 42448 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_383
timestamp 1698175906
transform 1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_387
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_403
timestamp 1698175906
transform 1 0 46480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_407
timestamp 1698175906
transform 1 0 46928 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_440
timestamp 1698175906
transform 1 0 50624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_448
timestamp 1698175906
transform 1 0 51520 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_452
timestamp 1698175906
transform 1 0 51968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698175906
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_457
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_88
timestamp 1698175906
transform 1 0 11200 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_92
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_94
timestamp 1698175906
transform 1 0 11872 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_97
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_107
timestamp 1698175906
transform 1 0 13328 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_123
timestamp 1698175906
transform 1 0 15120 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_131
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_135
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_174
timestamp 1698175906
transform 1 0 20832 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_190
timestamp 1698175906
transform 1 0 22624 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_194
timestamp 1698175906
transform 1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_202
timestamp 1698175906
transform 1 0 23968 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_224
timestamp 1698175906
transform 1 0 26432 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_240
timestamp 1698175906
transform 1 0 28224 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_256
timestamp 1698175906
transform 1 0 30016 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_264
timestamp 1698175906
transform 1 0 30912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698175906
transform 1 0 32368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698175906
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_288
timestamp 1698175906
transform 1 0 33600 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_296
timestamp 1698175906
transform 1 0 34496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_300
timestamp 1698175906
transform 1 0 34944 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_319
timestamp 1698175906
transform 1 0 37072 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_333
timestamp 1698175906
transform 1 0 38640 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698175906
transform 1 0 40432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_360
timestamp 1698175906
transform 1 0 41664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_362
timestamp 1698175906
transform 1 0 41888 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_368
timestamp 1698175906
transform 1 0 42560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_372
timestamp 1698175906
transform 1 0 43008 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_376
timestamp 1698175906
transform 1 0 43456 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_378
timestamp 1698175906
transform 1 0 43680 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_381
timestamp 1698175906
transform 1 0 44016 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_400
timestamp 1698175906
transform 1 0 46144 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698175906
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_422
timestamp 1698175906
transform 1 0 48608 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_438
timestamp 1698175906
transform 1 0 50400 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_446
timestamp 1698175906
transform 1 0 51296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_450
timestamp 1698175906
transform 1 0 51744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_452
timestamp 1698175906
transform 1 0 51968 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_461
timestamp 1698175906
transform 1 0 52976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_41
timestamp 1698175906
transform 1 0 5936 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_73
timestamp 1698175906
transform 1 0 9520 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_77
timestamp 1698175906
transform 1 0 9968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_79
timestamp 1698175906
transform 1 0 10192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_82
timestamp 1698175906
transform 1 0 10528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_84
timestamp 1698175906
transform 1 0 10752 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_119
timestamp 1698175906
transform 1 0 14672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_123
timestamp 1698175906
transform 1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_127
timestamp 1698175906
transform 1 0 15568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_131
timestamp 1698175906
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_164
timestamp 1698175906
transform 1 0 19712 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698175906
transform 1 0 20608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698175906
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_193
timestamp 1698175906
transform 1 0 22960 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_195
timestamp 1698175906
transform 1 0 23184 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_201
timestamp 1698175906
transform 1 0 23856 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_217
timestamp 1698175906
transform 1 0 25648 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_225
timestamp 1698175906
transform 1 0 26544 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_234
timestamp 1698175906
transform 1 0 27552 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_242
timestamp 1698175906
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698175906
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_253
timestamp 1698175906
transform 1 0 29680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_257
timestamp 1698175906
transform 1 0 30128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_273
timestamp 1698175906
transform 1 0 31920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_281
timestamp 1698175906
transform 1 0 32816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_285
timestamp 1698175906
transform 1 0 33264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_293
timestamp 1698175906
transform 1 0 34160 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_301
timestamp 1698175906
transform 1 0 35056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_305
timestamp 1698175906
transform 1 0 35504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_307
timestamp 1698175906
transform 1 0 35728 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698175906
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698175906
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_340
timestamp 1698175906
transform 1 0 39424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_379
timestamp 1698175906
transform 1 0 43792 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_383
timestamp 1698175906
transform 1 0 44240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_422
timestamp 1698175906
transform 1 0 48608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_426
timestamp 1698175906
transform 1 0 49056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_428
timestamp 1698175906
transform 1 0 49280 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_441
timestamp 1698175906
transform 1 0 50736 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_449
timestamp 1698175906
transform 1 0 51632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_453
timestamp 1698175906
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_457
timestamp 1698175906
transform 1 0 52528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_34
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_36
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_52
timestamp 1698175906
transform 1 0 7168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_56
timestamp 1698175906
transform 1 0 7616 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_64
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_85
timestamp 1698175906
transform 1 0 10864 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_92
timestamp 1698175906
transform 1 0 11648 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_146
timestamp 1698175906
transform 1 0 17696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_158
timestamp 1698175906
transform 1 0 19040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_162
timestamp 1698175906
transform 1 0 19488 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_194
timestamp 1698175906
transform 1 0 23072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_218
timestamp 1698175906
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_222
timestamp 1698175906
transform 1 0 26208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_261
timestamp 1698175906
transform 1 0 30576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_265
timestamp 1698175906
transform 1 0 31024 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_269
timestamp 1698175906
transform 1 0 31472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_298
timestamp 1698175906
transform 1 0 34720 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_302
timestamp 1698175906
transform 1 0 35168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_318
timestamp 1698175906
transform 1 0 36960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_322
timestamp 1698175906
transform 1 0 37408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_330
timestamp 1698175906
transform 1 0 38304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_344
timestamp 1698175906
transform 1 0 39872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_354
timestamp 1698175906
transform 1 0 40992 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_366
timestamp 1698175906
transform 1 0 42336 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_368
timestamp 1698175906
transform 1 0 42560 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_383
timestamp 1698175906
transform 1 0 44240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_385
timestamp 1698175906
transform 1 0 44464 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_400
timestamp 1698175906
transform 1 0 46144 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698175906
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_422
timestamp 1698175906
transform 1 0 48608 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_31
timestamp 1698175906
transform 1 0 4816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_48
timestamp 1698175906
transform 1 0 6720 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_64
timestamp 1698175906
transform 1 0 8512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_76
timestamp 1698175906
transform 1 0 9856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_80
timestamp 1698175906
transform 1 0 10304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_92
timestamp 1698175906
transform 1 0 11648 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_96
timestamp 1698175906
transform 1 0 12096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_98
timestamp 1698175906
transform 1 0 12320 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_117
timestamp 1698175906
transform 1 0 14448 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_144
timestamp 1698175906
transform 1 0 17472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_148
timestamp 1698175906
transform 1 0 17920 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_164
timestamp 1698175906
transform 1 0 19712 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_168
timestamp 1698175906
transform 1 0 20160 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_181
timestamp 1698175906
transform 1 0 21616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_189
timestamp 1698175906
transform 1 0 22512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_198
timestamp 1698175906
transform 1 0 23520 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_202
timestamp 1698175906
transform 1 0 23968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_204
timestamp 1698175906
transform 1 0 24192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_207
timestamp 1698175906
transform 1 0 24528 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_215
timestamp 1698175906
transform 1 0 25424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_217
timestamp 1698175906
transform 1 0 25648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_234
timestamp 1698175906
transform 1 0 27552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_238
timestamp 1698175906
transform 1 0 28000 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698175906
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698175906
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_253
timestamp 1698175906
transform 1 0 29680 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_261
timestamp 1698175906
transform 1 0 30576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_263
timestamp 1698175906
transform 1 0 30800 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_283
timestamp 1698175906
transform 1 0 33040 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_349
timestamp 1698175906
transform 1 0 40432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_368
timestamp 1698175906
transform 1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_372
timestamp 1698175906
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_376
timestamp 1698175906
transform 1 0 43456 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698175906
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_389
timestamp 1698175906
transform 1 0 44912 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_428
timestamp 1698175906
transform 1 0 49280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_432
timestamp 1698175906
transform 1 0 49728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_436
timestamp 1698175906
transform 1 0 50176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_438
timestamp 1698175906
transform 1 0 50400 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_443
timestamp 1698175906
transform 1 0 50960 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_451
timestamp 1698175906
transform 1 0 51856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_457
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698175906
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_26
timestamp 1698175906
transform 1 0 4256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_30
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_32
timestamp 1698175906
transform 1 0 4928 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_39
timestamp 1698175906
transform 1 0 5712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_61
timestamp 1698175906
transform 1 0 8176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_65
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698175906
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_104
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_118
timestamp 1698175906
transform 1 0 14560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_152
timestamp 1698175906
transform 1 0 18368 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_160
timestamp 1698175906
transform 1 0 19264 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_164
timestamp 1698175906
transform 1 0 19712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_173
timestamp 1698175906
transform 1 0 20720 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_189
timestamp 1698175906
transform 1 0 22512 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_238
timestamp 1698175906
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_242
timestamp 1698175906
transform 1 0 28448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_258
timestamp 1698175906
transform 1 0 30240 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_266
timestamp 1698175906
transform 1 0 31136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_305
timestamp 1698175906
transform 1 0 35504 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_315
timestamp 1698175906
transform 1 0 36624 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_323
timestamp 1698175906
transform 1 0 37520 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_338
timestamp 1698175906
transform 1 0 39200 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_392
timestamp 1698175906
transform 1 0 45248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_396
timestamp 1698175906
transform 1 0 45696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_398
timestamp 1698175906
transform 1 0 45920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_401
timestamp 1698175906
transform 1 0 46256 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_417
timestamp 1698175906
transform 1 0 48048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698175906
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_422
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_426
timestamp 1698175906
transform 1 0 49056 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_435
timestamp 1698175906
transform 1 0 50064 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_6
timestamp 1698175906
transform 1 0 2016 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_13
timestamp 1698175906
transform 1 0 2800 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_29
timestamp 1698175906
transform 1 0 4592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_33
timestamp 1698175906
transform 1 0 5040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_53
timestamp 1698175906
transform 1 0 7280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_66
timestamp 1698175906
transform 1 0 8736 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_82
timestamp 1698175906
transform 1 0 10528 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_85
timestamp 1698175906
transform 1 0 10864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_93
timestamp 1698175906
transform 1 0 11760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_95
timestamp 1698175906
transform 1 0 11984 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_98
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_102
timestamp 1698175906
transform 1 0 12768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698175906
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_113
timestamp 1698175906
transform 1 0 14000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_117
timestamp 1698175906
transform 1 0 14448 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_120
timestamp 1698175906
transform 1 0 14784 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_124
timestamp 1698175906
transform 1 0 15232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_136
timestamp 1698175906
transform 1 0 16576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_156
timestamp 1698175906
transform 1 0 18816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_160
timestamp 1698175906
transform 1 0 19264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_168
timestamp 1698175906
transform 1 0 20160 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698175906
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_193
timestamp 1698175906
transform 1 0 22960 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_228
timestamp 1698175906
transform 1 0 26880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_232
timestamp 1698175906
transform 1 0 27328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698175906
transform 1 0 28224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_255
timestamp 1698175906
transform 1 0 29904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_259
timestamp 1698175906
transform 1 0 30352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_290
timestamp 1698175906
transform 1 0 33824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_292
timestamp 1698175906
transform 1 0 34048 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_299
timestamp 1698175906
transform 1 0 34832 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698175906
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_321
timestamp 1698175906
transform 1 0 37296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_343
timestamp 1698175906
transform 1 0 39760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_347
timestamp 1698175906
transform 1 0 40208 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_357
timestamp 1698175906
transform 1 0 41328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_361
timestamp 1698175906
transform 1 0 41776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_363
timestamp 1698175906
transform 1 0 42000 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_370
timestamp 1698175906
transform 1 0 42784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_374
timestamp 1698175906
transform 1 0 43232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_382
timestamp 1698175906
transform 1 0 44128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698175906
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698175906
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_43
timestamp 1698175906
transform 1 0 6160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_51
timestamp 1698175906
transform 1 0 7056 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_76
timestamp 1698175906
transform 1 0 9856 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_83
timestamp 1698175906
transform 1 0 10640 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_96
timestamp 1698175906
transform 1 0 12096 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_103
timestamp 1698175906
transform 1 0 12880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_107
timestamp 1698175906
transform 1 0 13328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_139
timestamp 1698175906
transform 1 0 16912 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_158
timestamp 1698175906
transform 1 0 19040 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_166
timestamp 1698175906
transform 1 0 19936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_170
timestamp 1698175906
transform 1 0 20384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_172
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_177
timestamp 1698175906
transform 1 0 21168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_253
timestamp 1698175906
transform 1 0 29680 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_269
timestamp 1698175906
transform 1 0 31472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698175906
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_298
timestamp 1698175906
transform 1 0 34720 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_302
timestamp 1698175906
transform 1 0 35168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_304
timestamp 1698175906
transform 1 0 35392 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_317
timestamp 1698175906
transform 1 0 36848 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_325
timestamp 1698175906
transform 1 0 37744 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_329
timestamp 1698175906
transform 1 0 38192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_352
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_389
timestamp 1698175906
transform 1 0 44912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_393
timestamp 1698175906
transform 1 0 45360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_407
timestamp 1698175906
transform 1 0 46928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_415
timestamp 1698175906
transform 1 0 47824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698175906
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_422
timestamp 1698175906
transform 1 0 48608 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_454
timestamp 1698175906
transform 1 0 52192 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_462
timestamp 1698175906
transform 1 0 53088 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_41
timestamp 1698175906
transform 1 0 5936 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_50
timestamp 1698175906
transform 1 0 6944 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_58
timestamp 1698175906
transform 1 0 7840 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_72
timestamp 1698175906
transform 1 0 9408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_76
timestamp 1698175906
transform 1 0 9856 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_92
timestamp 1698175906
transform 1 0 11648 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_100
timestamp 1698175906
transform 1 0 12544 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_104
timestamp 1698175906
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 14224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_119
timestamp 1698175906
transform 1 0 14672 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_133
timestamp 1698175906
transform 1 0 16240 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698175906
transform 1 0 16688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698175906
transform 1 0 16912 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_156
timestamp 1698175906
transform 1 0 18816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_160
timestamp 1698175906
transform 1 0 19264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_168
timestamp 1698175906
transform 1 0 20160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_193
timestamp 1698175906
transform 1 0 22960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_201
timestamp 1698175906
transform 1 0 23856 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_207
timestamp 1698175906
transform 1 0 24528 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_215
timestamp 1698175906
transform 1 0 25424 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_224
timestamp 1698175906
transform 1 0 26432 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 28224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_249
timestamp 1698175906
transform 1 0 29232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_252
timestamp 1698175906
transform 1 0 29568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_260
timestamp 1698175906
transform 1 0 30464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_264
timestamp 1698175906
transform 1 0 30912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_278
timestamp 1698175906
transform 1 0 32480 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_294
timestamp 1698175906
transform 1 0 34272 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_302
timestamp 1698175906
transform 1 0 35168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_306
timestamp 1698175906
transform 1 0 35616 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698175906
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698175906
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_325
timestamp 1698175906
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_359
timestamp 1698175906
transform 1 0 41552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_367
timestamp 1698175906
transform 1 0 42448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_371
timestamp 1698175906
transform 1 0 42896 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_379
timestamp 1698175906
transform 1 0 43792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_383
timestamp 1698175906
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_409
timestamp 1698175906
transform 1 0 47152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_413
timestamp 1698175906
transform 1 0 47600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_415
timestamp 1698175906
transform 1 0 47824 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_445
timestamp 1698175906
transform 1 0 51184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_449
timestamp 1698175906
transform 1 0 51632 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_453
timestamp 1698175906
transform 1 0 52080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_34
timestamp 1698175906
transform 1 0 5152 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_38
timestamp 1698175906
transform 1 0 5600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_45
timestamp 1698175906
transform 1 0 6384 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_67
timestamp 1698175906
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698175906
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_76
timestamp 1698175906
transform 1 0 9856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_78
timestamp 1698175906
transform 1 0 10080 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_89
timestamp 1698175906
transform 1 0 11312 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_105
timestamp 1698175906
transform 1 0 13104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_107
timestamp 1698175906
transform 1 0 13328 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_152
timestamp 1698175906
transform 1 0 18368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_183
timestamp 1698175906
transform 1 0 21840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_187
timestamp 1698175906
transform 1 0 22288 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_203
timestamp 1698175906
transform 1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_228
timestamp 1698175906
transform 1 0 26880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_236
timestamp 1698175906
transform 1 0 27776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_240
timestamp 1698175906
transform 1 0 28224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_250
timestamp 1698175906
transform 1 0 29344 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_284
timestamp 1698175906
transform 1 0 33152 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_289
timestamp 1698175906
transform 1 0 33712 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_296
timestamp 1698175906
transform 1 0 34496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_300
timestamp 1698175906
transform 1 0 34944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_344
timestamp 1698175906
transform 1 0 39872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698175906
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_385
timestamp 1698175906
transform 1 0 44464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_389
timestamp 1698175906
transform 1 0 44912 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_405
timestamp 1698175906
transform 1 0 46704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_413
timestamp 1698175906
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_417
timestamp 1698175906
transform 1 0 48048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698175906
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_428
timestamp 1698175906
transform 1 0 49280 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_458
timestamp 1698175906
transform 1 0 52640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_462
timestamp 1698175906
transform 1 0 53088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_464
timestamp 1698175906
transform 1 0 53312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_18
timestamp 1698175906
transform 1 0 3360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_22
timestamp 1698175906
transform 1 0 3808 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_51
timestamp 1698175906
transform 1 0 7056 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_67
timestamp 1698175906
transform 1 0 8848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_71
timestamp 1698175906
transform 1 0 9296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_111
timestamp 1698175906
transform 1 0 13776 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_119
timestamp 1698175906
transform 1 0 14672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_123
timestamp 1698175906
transform 1 0 15120 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_130
timestamp 1698175906
transform 1 0 15904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_138
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_140
timestamp 1698175906
transform 1 0 17024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_147
timestamp 1698175906
transform 1 0 17808 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_163
timestamp 1698175906
transform 1 0 19600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698175906
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698175906
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698175906
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_200
timestamp 1698175906
transform 1 0 23744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_210
timestamp 1698175906
transform 1 0 24864 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_219
timestamp 1698175906
transform 1 0 25872 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_235
timestamp 1698175906
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_279
timestamp 1698175906
transform 1 0 32592 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_295
timestamp 1698175906
transform 1 0 34384 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_308
timestamp 1698175906
transform 1 0 35840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698175906
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698175906
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_321
timestamp 1698175906
transform 1 0 37296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698175906
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_391
timestamp 1698175906
transform 1 0 45136 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_407
timestamp 1698175906
transform 1 0 46928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_415
timestamp 1698175906
transform 1 0 47824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_419
timestamp 1698175906
transform 1 0 48272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_429
timestamp 1698175906
transform 1 0 49392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_443
timestamp 1698175906
transform 1 0 50960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_447
timestamp 1698175906
transform 1 0 51408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_449
timestamp 1698175906
transform 1 0 51632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_31
timestamp 1698175906
transform 1 0 4816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_35
timestamp 1698175906
transform 1 0 5264 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_53
timestamp 1698175906
transform 1 0 7280 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_57
timestamp 1698175906
transform 1 0 7728 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_65
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698175906
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_114
timestamp 1698175906
transform 1 0 14112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_126
timestamp 1698175906
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_152
timestamp 1698175906
transform 1 0 18368 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_160
timestamp 1698175906
transform 1 0 19264 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_164
timestamp 1698175906
transform 1 0 19712 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_170
timestamp 1698175906
transform 1 0 20384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_172
timestamp 1698175906
transform 1 0 20608 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 24528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_241
timestamp 1698175906
transform 1 0 28336 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_273
timestamp 1698175906
transform 1 0 31920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_275
timestamp 1698175906
transform 1 0 32144 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_298
timestamp 1698175906
transform 1 0 34720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_306
timestamp 1698175906
transform 1 0 35616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_310
timestamp 1698175906
transform 1 0 36064 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_315
timestamp 1698175906
transform 1 0 36624 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_323
timestamp 1698175906
transform 1 0 37520 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_329
timestamp 1698175906
transform 1 0 38192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698175906
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_380
timestamp 1698175906
transform 1 0 43904 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_392
timestamp 1698175906
transform 1 0 45248 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_408
timestamp 1698175906
transform 1 0 47040 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698175906
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_431
timestamp 1698175906
transform 1 0 49616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_439
timestamp 1698175906
transform 1 0 50512 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_443
timestamp 1698175906
transform 1 0 50960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_445
timestamp 1698175906
transform 1 0 51184 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_448
timestamp 1698175906
transform 1 0 51520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_452
timestamp 1698175906
transform 1 0 51968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_456
timestamp 1698175906
transform 1 0 52416 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_56
timestamp 1698175906
transform 1 0 7616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_60
timestamp 1698175906
transform 1 0 8064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_67
timestamp 1698175906
transform 1 0 8848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_71
timestamp 1698175906
transform 1 0 9296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_81
timestamp 1698175906
transform 1 0 10416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_85
timestamp 1698175906
transform 1 0 10864 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_139
timestamp 1698175906
transform 1 0 16912 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_142
timestamp 1698175906
transform 1 0 17248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_209
timestamp 1698175906
transform 1 0 24752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_212
timestamp 1698175906
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_214
timestamp 1698175906
transform 1 0 25312 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_220
timestamp 1698175906
transform 1 0 25984 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_236
timestamp 1698175906
transform 1 0 27776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_240
timestamp 1698175906
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_242
timestamp 1698175906
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_282
timestamp 1698175906
transform 1 0 32928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_286
timestamp 1698175906
transform 1 0 33376 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_297
timestamp 1698175906
transform 1 0 34608 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_325
timestamp 1698175906
transform 1 0 37744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_327
timestamp 1698175906
transform 1 0 37968 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_330
timestamp 1698175906
transform 1 0 38304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698175906
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_391
timestamp 1698175906
transform 1 0 45136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_395
timestamp 1698175906
transform 1 0 45584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_425
timestamp 1698175906
transform 1 0 48944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_429
timestamp 1698175906
transform 1 0 49392 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_437
timestamp 1698175906
transform 1 0 50288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_453
timestamp 1698175906
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_457
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_34
timestamp 1698175906
transform 1 0 5152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_38
timestamp 1698175906
transform 1 0 5600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_40
timestamp 1698175906
transform 1 0 5824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_56
timestamp 1698175906
transform 1 0 7616 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_76
timestamp 1698175906
transform 1 0 9856 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_92
timestamp 1698175906
transform 1 0 11648 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_96
timestamp 1698175906
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_131
timestamp 1698175906
transform 1 0 16016 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_216
timestamp 1698175906
transform 1 0 25536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_224
timestamp 1698175906
transform 1 0 26432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_235
timestamp 1698175906
transform 1 0 27664 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_251
timestamp 1698175906
transform 1 0 29456 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_259
timestamp 1698175906
transform 1 0 30352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_263
timestamp 1698175906
transform 1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_313
timestamp 1698175906
transform 1 0 36400 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_333
timestamp 1698175906
transform 1 0 38640 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698175906
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1698175906
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_381
timestamp 1698175906
transform 1 0 44016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_393
timestamp 1698175906
transform 1 0 45360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_401
timestamp 1698175906
transform 1 0 46256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_409
timestamp 1698175906
transform 1 0 47152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_413
timestamp 1698175906
transform 1 0 47600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_417
timestamp 1698175906
transform 1 0 48048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698175906
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_422
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_426
timestamp 1698175906
transform 1 0 49056 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_433
timestamp 1698175906
transform 1 0 49840 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_437
timestamp 1698175906
transform 1 0 50288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_439
timestamp 1698175906
transform 1 0 50512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_462
timestamp 1698175906
transform 1 0 53088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_464
timestamp 1698175906
transform 1 0 53312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_31
timestamp 1698175906
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_53
timestamp 1698175906
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_61
timestamp 1698175906
transform 1 0 8176 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_68
timestamp 1698175906
transform 1 0 8960 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_84
timestamp 1698175906
transform 1 0 10752 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_88
timestamp 1698175906
transform 1 0 11200 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_95
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_139
timestamp 1698175906
transform 1 0 16912 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_142
timestamp 1698175906
transform 1 0 17248 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_158
timestamp 1698175906
transform 1 0 19040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_166
timestamp 1698175906
transform 1 0 19936 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_207
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_252
timestamp 1698175906
transform 1 0 29568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_256
timestamp 1698175906
transform 1 0 30016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_260
timestamp 1698175906
transform 1 0 30464 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_276
timestamp 1698175906
transform 1 0 32256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_282
timestamp 1698175906
transform 1 0 32928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_286
timestamp 1698175906
transform 1 0 33376 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_292
timestamp 1698175906
transform 1 0 34048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_296
timestamp 1698175906
transform 1 0 34496 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_329
timestamp 1698175906
transform 1 0 38192 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_333
timestamp 1698175906
transform 1 0 38640 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_336
timestamp 1698175906
transform 1 0 38976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_377
timestamp 1698175906
transform 1 0 43568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_381
timestamp 1698175906
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_391
timestamp 1698175906
transform 1 0 45136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_395
timestamp 1698175906
transform 1 0 45584 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_403
timestamp 1698175906
transform 1 0 46480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_409
timestamp 1698175906
transform 1 0 47152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_416
timestamp 1698175906
transform 1 0 47936 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_443
timestamp 1698175906
transform 1 0 50960 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_451
timestamp 1698175906
transform 1 0 51856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_457
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_10
timestamp 1698175906
transform 1 0 2464 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_17
timestamp 1698175906
transform 1 0 3248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_21
timestamp 1698175906
transform 1 0 3696 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_29
timestamp 1698175906
transform 1 0 4592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_33
timestamp 1698175906
transform 1 0 5040 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_42
timestamp 1698175906
transform 1 0 6048 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_63
timestamp 1698175906
transform 1 0 8400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698175906
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698175906
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_88
timestamp 1698175906
transform 1 0 11200 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 12992 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_112
timestamp 1698175906
transform 1 0 13888 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_116
timestamp 1698175906
transform 1 0 14336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_130
timestamp 1698175906
transform 1 0 15904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_205
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_220
timestamp 1698175906
transform 1 0 25984 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_229
timestamp 1698175906
transform 1 0 26992 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_245
timestamp 1698175906
transform 1 0 28784 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_253
timestamp 1698175906
transform 1 0 29680 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_255
timestamp 1698175906
transform 1 0 29904 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_262
timestamp 1698175906
transform 1 0 30688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_266
timestamp 1698175906
transform 1 0 31136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_270
timestamp 1698175906
transform 1 0 31584 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_288
timestamp 1698175906
transform 1 0 33600 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_304
timestamp 1698175906
transform 1 0 35392 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_312
timestamp 1698175906
transform 1 0 36288 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_316
timestamp 1698175906
transform 1 0 36736 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_323
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_327
timestamp 1698175906
transform 1 0 37968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_335
timestamp 1698175906
transform 1 0 38864 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_339
timestamp 1698175906
transform 1 0 39312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_341
timestamp 1698175906
transform 1 0 39536 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_368
timestamp 1698175906
transform 1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_372
timestamp 1698175906
transform 1 0 43008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_374
timestamp 1698175906
transform 1 0 43232 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_397
timestamp 1698175906
transform 1 0 45808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698175906
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_434
timestamp 1698175906
transform 1 0 49952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_49
timestamp 1698175906
transform 1 0 6832 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_65
timestamp 1698175906
transform 1 0 8624 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_73
timestamp 1698175906
transform 1 0 9520 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_123
timestamp 1698175906
transform 1 0 15120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_131
timestamp 1698175906
transform 1 0 16016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_141
timestamp 1698175906
transform 1 0 17136 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_193
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_202
timestamp 1698175906
transform 1 0 23968 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_234
timestamp 1698175906
transform 1 0 27552 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_242
timestamp 1698175906
transform 1 0 28448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_252
timestamp 1698175906
transform 1 0 29568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_290
timestamp 1698175906
transform 1 0 33824 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_294
timestamp 1698175906
transform 1 0 34272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_301
timestamp 1698175906
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_319
timestamp 1698175906
transform 1 0 37072 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_374
timestamp 1698175906
transform 1 0 43232 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_378
timestamp 1698175906
transform 1 0 43680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_382
timestamp 1698175906
transform 1 0 44128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698175906
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_387
timestamp 1698175906
transform 1 0 44688 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_396
timestamp 1698175906
transform 1 0 45696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_400
timestamp 1698175906
transform 1 0 46144 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_416
timestamp 1698175906
transform 1 0 47936 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_424
timestamp 1698175906
transform 1 0 48832 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_428
timestamp 1698175906
transform 1 0 49280 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_435
timestamp 1698175906
transform 1 0 50064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_439
timestamp 1698175906
transform 1 0 50512 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_457
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_16
timestamp 1698175906
transform 1 0 3136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_20
timestamp 1698175906
transform 1 0 3584 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_30
timestamp 1698175906
transform 1 0 4704 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_33
timestamp 1698175906
transform 1 0 5040 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_56
timestamp 1698175906
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_64
timestamp 1698175906
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_76
timestamp 1698175906
transform 1 0 9856 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_92
timestamp 1698175906
transform 1 0 11648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_100
timestamp 1698175906
transform 1 0 12544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_104
timestamp 1698175906
transform 1 0 12992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_106
timestamp 1698175906
transform 1 0 13216 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_144
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_153
timestamp 1698175906
transform 1 0 18480 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_169
timestamp 1698175906
transform 1 0 20272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_204
timestamp 1698175906
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_220
timestamp 1698175906
transform 1 0 25984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_224
timestamp 1698175906
transform 1 0 26432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_231
timestamp 1698175906
transform 1 0 27216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_235
timestamp 1698175906
transform 1 0 27664 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_251
timestamp 1698175906
transform 1 0 29456 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_259
timestamp 1698175906
transform 1 0 30352 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_261
timestamp 1698175906
transform 1 0 30576 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_264
timestamp 1698175906
transform 1 0 30912 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_290
timestamp 1698175906
transform 1 0 33824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_292
timestamp 1698175906
transform 1 0 34048 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_388
timestamp 1698175906
transform 1 0 44800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_392
timestamp 1698175906
transform 1 0 45248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_408
timestamp 1698175906
transform 1 0 47040 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_412
timestamp 1698175906
transform 1 0 47488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698175906
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_430
timestamp 1698175906
transform 1 0 49504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_440
timestamp 1698175906
transform 1 0 50624 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_456
timestamp 1698175906
transform 1 0 52416 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698175906
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_46
timestamp 1698175906
transform 1 0 6496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_50
timestamp 1698175906
transform 1 0 6944 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_86
timestamp 1698175906
transform 1 0 10976 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_102
timestamp 1698175906
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698175906
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_118
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_122
timestamp 1698175906
transform 1 0 15008 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_126
timestamp 1698175906
transform 1 0 15456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_133
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_141
timestamp 1698175906
transform 1 0 17136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_193
timestamp 1698175906
transform 1 0 22960 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_201
timestamp 1698175906
transform 1 0 23856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698175906
transform 1 0 28224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_257
timestamp 1698175906
transform 1 0 30128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_261
timestamp 1698175906
transform 1 0 30576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_302
timestamp 1698175906
transform 1 0 35168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_310
timestamp 1698175906
transform 1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_312
timestamp 1698175906
transform 1 0 36288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_319
timestamp 1698175906
transform 1 0 37072 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_369
timestamp 1698175906
transform 1 0 42672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_379
timestamp 1698175906
transform 1 0 43792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698175906
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_450
timestamp 1698175906
transform 1 0 51744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_452
timestamp 1698175906
transform 1 0 51968 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_463
timestamp 1698175906
transform 1 0 53200 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698175906
transform 1 0 3360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_26
timestamp 1698175906
transform 1 0 4256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_36
timestamp 1698175906
transform 1 0 5376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_40
timestamp 1698175906
transform 1 0 5824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_47
timestamp 1698175906
transform 1 0 6608 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_63
timestamp 1698175906
transform 1 0 8400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698175906
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698175906
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_76
timestamp 1698175906
transform 1 0 9856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_92
timestamp 1698175906
transform 1 0 11648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_106
timestamp 1698175906
transform 1 0 13216 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698175906
transform 1 0 19264 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_175
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_179
timestamp 1698175906
transform 1 0 21392 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_195
timestamp 1698175906
transform 1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698175906
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698175906
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_228
timestamp 1698175906
transform 1 0 26880 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_234
timestamp 1698175906
transform 1 0 27552 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_266
timestamp 1698175906
transform 1 0 31136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_272
timestamp 1698175906
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_316
timestamp 1698175906
transform 1 0 36736 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_323
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_327
timestamp 1698175906
transform 1 0 37968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_335
timestamp 1698175906
transform 1 0 38864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_337
timestamp 1698175906
transform 1 0 39088 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_344
timestamp 1698175906
transform 1 0 39872 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698175906
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_366
timestamp 1698175906
transform 1 0 42336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_370
timestamp 1698175906
transform 1 0 42784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_372
timestamp 1698175906
transform 1 0 43008 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_387
timestamp 1698175906
transform 1 0 44688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_391
timestamp 1698175906
transform 1 0 45136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_395
timestamp 1698175906
transform 1 0 45584 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_411
timestamp 1698175906
transform 1 0 47376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_415
timestamp 1698175906
transform 1 0 47824 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_418
timestamp 1698175906
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_435
timestamp 1698175906
transform 1 0 50064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_16
timestamp 1698175906
transform 1 0 3136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_20
timestamp 1698175906
transform 1 0 3584 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_43
timestamp 1698175906
transform 1 0 6160 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_51
timestamp 1698175906
transform 1 0 7056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_55
timestamp 1698175906
transform 1 0 7504 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_62
timestamp 1698175906
transform 1 0 8288 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_78
timestamp 1698175906
transform 1 0 10080 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_86
timestamp 1698175906
transform 1 0 10976 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_96
timestamp 1698175906
transform 1 0 12096 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698175906
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_140
timestamp 1698175906
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_144
timestamp 1698175906
transform 1 0 17472 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_160
timestamp 1698175906
transform 1 0 19264 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 20160 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 20608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698175906
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_218
timestamp 1698175906
transform 1 0 25760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_222
timestamp 1698175906
transform 1 0 26208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_232
timestamp 1698175906
transform 1 0 27328 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_240
timestamp 1698175906
transform 1 0 28224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_278
timestamp 1698175906
transform 1 0 32480 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_294
timestamp 1698175906
transform 1 0 34272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_296
timestamp 1698175906
transform 1 0 34496 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_302
timestamp 1698175906
transform 1 0 35168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_322
timestamp 1698175906
transform 1 0 37408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_330
timestamp 1698175906
transform 1 0 38304 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_336
timestamp 1698175906
transform 1 0 38976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_344
timestamp 1698175906
transform 1 0 39872 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_348
timestamp 1698175906
transform 1 0 40320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_375
timestamp 1698175906
transform 1 0 43344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_397
timestamp 1698175906
transform 1 0 45808 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_409
timestamp 1698175906
transform 1 0 47152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_417
timestamp 1698175906
transform 1 0 48048 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_420
timestamp 1698175906
transform 1 0 48384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_428
timestamp 1698175906
transform 1 0 49280 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_432
timestamp 1698175906
transform 1 0 49728 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_440
timestamp 1698175906
transform 1 0 50624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_444
timestamp 1698175906
transform 1 0 51072 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_452
timestamp 1698175906
transform 1 0 51968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_454
timestamp 1698175906
transform 1 0 52192 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_31
timestamp 1698175906
transform 1 0 4816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_43
timestamp 1698175906
transform 1 0 6160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_45
timestamp 1698175906
transform 1 0 6384 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_52
timestamp 1698175906
transform 1 0 7168 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_111
timestamp 1698175906
transform 1 0 13776 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_127
timestamp 1698175906
transform 1 0 15568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698175906
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_150
timestamp 1698175906
transform 1 0 18144 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_160
timestamp 1698175906
transform 1 0 19264 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_164
timestamp 1698175906
transform 1 0 19712 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_196
timestamp 1698175906
transform 1 0 23296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_200
timestamp 1698175906
transform 1 0 23744 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_230
timestamp 1698175906
transform 1 0 27104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_234
timestamp 1698175906
transform 1 0 27552 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_256
timestamp 1698175906
transform 1 0 30016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_260
timestamp 1698175906
transform 1 0 30464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_264
timestamp 1698175906
transform 1 0 30912 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698175906
transform 1 0 33824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_302
timestamp 1698175906
transform 1 0 35168 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_360
timestamp 1698175906
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_362
timestamp 1698175906
transform 1 0 41888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_385
timestamp 1698175906
transform 1 0 44464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_389
timestamp 1698175906
transform 1 0 44912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_427
timestamp 1698175906
transform 1 0 49168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_431
timestamp 1698175906
transform 1 0 49616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_435
timestamp 1698175906
transform 1 0 50064 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_443
timestamp 1698175906
transform 1 0 50960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_445
timestamp 1698175906
transform 1 0 51184 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_454
timestamp 1698175906
transform 1 0 52192 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_462
timestamp 1698175906
transform 1 0 53088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_52
timestamp 1698175906
transform 1 0 7168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_60
timestamp 1698175906
transform 1 0 8064 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_64
timestamp 1698175906
transform 1 0 8512 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_85
timestamp 1698175906
transform 1 0 10864 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_139
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_143
timestamp 1698175906
transform 1 0 17360 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_166
timestamp 1698175906
transform 1 0 19936 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_213
timestamp 1698175906
transform 1 0 25200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_215
timestamp 1698175906
transform 1 0 25424 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_230
timestamp 1698175906
transform 1 0 27104 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_253
timestamp 1698175906
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_257
timestamp 1698175906
transform 1 0 30128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_261
timestamp 1698175906
transform 1 0 30576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_296
timestamp 1698175906
transform 1 0 34496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_300
timestamp 1698175906
transform 1 0 34944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_304
timestamp 1698175906
transform 1 0 35392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698175906
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_349
timestamp 1698175906
transform 1 0 40432 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_365
timestamp 1698175906
transform 1 0 42224 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_373
timestamp 1698175906
transform 1 0 43120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_377
timestamp 1698175906
transform 1 0 43568 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_387
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_419
timestamp 1698175906
transform 1 0 48272 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_422
timestamp 1698175906
transform 1 0 48608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_426
timestamp 1698175906
transform 1 0 49056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698175906
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_34
timestamp 1698175906
transform 1 0 5152 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_44
timestamp 1698175906
transform 1 0 6272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_53
timestamp 1698175906
transform 1 0 7280 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698175906
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_78
timestamp 1698175906
transform 1 0 10080 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_86
timestamp 1698175906
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_105
timestamp 1698175906
transform 1 0 13104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_109
timestamp 1698175906
transform 1 0 13552 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_117
timestamp 1698175906
transform 1 0 14448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_121
timestamp 1698175906
transform 1 0 14896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_129
timestamp 1698175906
transform 1 0 15792 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698175906
transform 1 0 18592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_158
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_190
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_201
timestamp 1698175906
transform 1 0 23856 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_224
timestamp 1698175906
transform 1 0 26432 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_256
timestamp 1698175906
transform 1 0 30016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_260
timestamp 1698175906
transform 1 0 30464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_262
timestamp 1698175906
transform 1 0 30688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_332
timestamp 1698175906
transform 1 0 38528 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698175906
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_381
timestamp 1698175906
transform 1 0 44016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_393
timestamp 1698175906
transform 1 0 45360 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_409
timestamp 1698175906
transform 1 0 47152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_417
timestamp 1698175906
transform 1 0 48048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698175906
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_422
timestamp 1698175906
transform 1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_424
timestamp 1698175906
transform 1 0 48832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_430
timestamp 1698175906
transform 1 0 49504 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_436
timestamp 1698175906
transform 1 0 50176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_444
timestamp 1698175906
transform 1 0 51072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_453
timestamp 1698175906
transform 1 0 52080 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_461
timestamp 1698175906
transform 1 0 52976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_18
timestamp 1698175906
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_26
timestamp 1698175906
transform 1 0 4256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_30
timestamp 1698175906
transform 1 0 4704 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_33
timestamp 1698175906
transform 1 0 5040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_49
timestamp 1698175906
transform 1 0 6832 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_81
timestamp 1698175906
transform 1 0 10416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_85
timestamp 1698175906
transform 1 0 10864 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_136
timestamp 1698175906
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_140
timestamp 1698175906
transform 1 0 17024 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 20608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_191
timestamp 1698175906
transform 1 0 22736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_224
timestamp 1698175906
transform 1 0 26432 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_255
timestamp 1698175906
transform 1 0 29904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_274
timestamp 1698175906
transform 1 0 32032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_278
timestamp 1698175906
transform 1 0 32480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_282
timestamp 1698175906
transform 1 0 32928 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_290
timestamp 1698175906
transform 1 0 33824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_294
timestamp 1698175906
transform 1 0 34272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_310
timestamp 1698175906
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698175906
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_322
timestamp 1698175906
transform 1 0 37408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_341
timestamp 1698175906
transform 1 0 39536 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_343
timestamp 1698175906
transform 1 0 39760 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_352
timestamp 1698175906
transform 1 0 40768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_356
timestamp 1698175906
transform 1 0 41216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_360
timestamp 1698175906
transform 1 0 41664 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_376
timestamp 1698175906
transform 1 0 43456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_380
timestamp 1698175906
transform 1 0 43904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_382
timestamp 1698175906
transform 1 0 44128 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_395
timestamp 1698175906
transform 1 0 45584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_397
timestamp 1698175906
transform 1 0 45808 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_400
timestamp 1698175906
transform 1 0 46144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_402
timestamp 1698175906
transform 1 0 46368 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_415
timestamp 1698175906
transform 1 0 47824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_419
timestamp 1698175906
transform 1 0 48272 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698175906
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_37
timestamp 1698175906
transform 1 0 5488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_59
timestamp 1698175906
transform 1 0 7952 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_63
timestamp 1698175906
transform 1 0 8400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698175906
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698175906
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_76
timestamp 1698175906
transform 1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_78
timestamp 1698175906
transform 1 0 10080 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_85
timestamp 1698175906
transform 1 0 10864 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_117
timestamp 1698175906
transform 1 0 14448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_133
timestamp 1698175906
transform 1 0 16240 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_137
timestamp 1698175906
transform 1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698175906
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698175906
transform 1 0 18144 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_166
timestamp 1698175906
transform 1 0 19936 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_170
timestamp 1698175906
transform 1 0 20384 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_178
timestamp 1698175906
transform 1 0 21280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_185
timestamp 1698175906
transform 1 0 22064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_189
timestamp 1698175906
transform 1 0 22512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_290
timestamp 1698175906
transform 1 0 33824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_303
timestamp 1698175906
transform 1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_307
timestamp 1698175906
transform 1 0 35728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_311
timestamp 1698175906
transform 1 0 36176 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_317
timestamp 1698175906
transform 1 0 36848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_333
timestamp 1698175906
transform 1 0 38640 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_341
timestamp 1698175906
transform 1 0 39536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_356
timestamp 1698175906
transform 1 0 41216 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_372
timestamp 1698175906
transform 1 0 43008 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_380
timestamp 1698175906
transform 1 0 43904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_382
timestamp 1698175906
transform 1 0 44128 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_398
timestamp 1698175906
transform 1 0 45920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_400
timestamp 1698175906
transform 1 0 46144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_406
timestamp 1698175906
transform 1 0 46816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_410
timestamp 1698175906
transform 1 0 47264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_412
timestamp 1698175906
transform 1 0 47488 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_415
timestamp 1698175906
transform 1 0 47824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698175906
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_422
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_424
timestamp 1698175906
transform 1 0 48832 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_427
timestamp 1698175906
transform 1 0 49168 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_431
timestamp 1698175906
transform 1 0 49616 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_433
timestamp 1698175906
transform 1 0 49840 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_47
timestamp 1698175906
transform 1 0 6608 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_55
timestamp 1698175906
transform 1 0 7504 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_59
timestamp 1698175906
transform 1 0 7952 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_70
timestamp 1698175906
transform 1 0 9184 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_74
timestamp 1698175906
transform 1 0 9632 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_76
timestamp 1698175906
transform 1 0 9856 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_81
timestamp 1698175906
transform 1 0 10416 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_111
timestamp 1698175906
transform 1 0 13776 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_127
timestamp 1698175906
transform 1 0 15568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_137
timestamp 1698175906
transform 1 0 16688 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_153
timestamp 1698175906
transform 1 0 18480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_157
timestamp 1698175906
transform 1 0 18928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698175906
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_187
timestamp 1698175906
transform 1 0 22288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_193
timestamp 1698175906
transform 1 0 22960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_197
timestamp 1698175906
transform 1 0 23408 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_213
timestamp 1698175906
transform 1 0 25200 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_221
timestamp 1698175906
transform 1 0 26096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_225
timestamp 1698175906
transform 1 0 26544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_227
timestamp 1698175906
transform 1 0 26768 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_236
timestamp 1698175906
transform 1 0 27776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_240
timestamp 1698175906
transform 1 0 28224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_255
timestamp 1698175906
transform 1 0 29904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_259
timestamp 1698175906
transform 1 0 30352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_298
timestamp 1698175906
transform 1 0 34720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_302
timestamp 1698175906
transform 1 0 35168 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_306
timestamp 1698175906
transform 1 0 35616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_330
timestamp 1698175906
transform 1 0 38304 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_334
timestamp 1698175906
transform 1 0 38752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_343
timestamp 1698175906
transform 1 0 39760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_355
timestamp 1698175906
transform 1 0 41104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_359
timestamp 1698175906
transform 1 0 41552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_363
timestamp 1698175906
transform 1 0 42000 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_379
timestamp 1698175906
transform 1 0 43792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698175906
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_387
timestamp 1698175906
transform 1 0 44688 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_395
timestamp 1698175906
transform 1 0 45584 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_414
timestamp 1698175906
transform 1 0 47712 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_433
timestamp 1698175906
transform 1 0 49840 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_449
timestamp 1698175906
transform 1 0 51632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_453
timestamp 1698175906
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_457
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_34
timestamp 1698175906
transform 1 0 5152 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_38
timestamp 1698175906
transform 1 0 5600 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_52
timestamp 1698175906
transform 1 0 7168 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_60
timestamp 1698175906
transform 1 0 8064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_88
timestamp 1698175906
transform 1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_92
timestamp 1698175906
transform 1 0 11648 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_99
timestamp 1698175906
transform 1 0 12432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_135
timestamp 1698175906
transform 1 0 16464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_137
timestamp 1698175906
transform 1 0 16688 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_172
timestamp 1698175906
transform 1 0 20608 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_204
timestamp 1698175906
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698175906
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698175906
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_242
timestamp 1698175906
transform 1 0 28448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_244
timestamp 1698175906
transform 1 0 28672 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_247
timestamp 1698175906
transform 1 0 29008 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_255
timestamp 1698175906
transform 1 0 29904 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_259
timestamp 1698175906
transform 1 0 30352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_273
timestamp 1698175906
transform 1 0 31920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698175906
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698175906
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_290
timestamp 1698175906
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_303
timestamp 1698175906
transform 1 0 35280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_336
timestamp 1698175906
transform 1 0 38976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_340
timestamp 1698175906
transform 1 0 39424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_360
timestamp 1698175906
transform 1 0 41664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_392
timestamp 1698175906
transform 1 0 45248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_396
timestamp 1698175906
transform 1 0 45696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_400
timestamp 1698175906
transform 1 0 46144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_402
timestamp 1698175906
transform 1 0 46368 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_413
timestamp 1698175906
transform 1 0 47600 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_422
timestamp 1698175906
transform 1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_424
timestamp 1698175906
transform 1 0 48832 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_454
timestamp 1698175906
transform 1 0 52192 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_458
timestamp 1698175906
transform 1 0 52640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_462
timestamp 1698175906
transform 1 0 53088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_31
timestamp 1698175906
transform 1 0 4816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_41
timestamp 1698175906
transform 1 0 5936 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_50
timestamp 1698175906
transform 1 0 6944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_54
timestamp 1698175906
transform 1 0 7392 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_77
timestamp 1698175906
transform 1 0 9968 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_93
timestamp 1698175906
transform 1 0 11760 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_115
timestamp 1698175906
transform 1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_119
timestamp 1698175906
transform 1 0 14672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_121
timestamp 1698175906
transform 1 0 14896 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_134
timestamp 1698175906
transform 1 0 16352 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_140
timestamp 1698175906
transform 1 0 17024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_144
timestamp 1698175906
transform 1 0 17472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_158
timestamp 1698175906
transform 1 0 19040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_162
timestamp 1698175906
transform 1 0 19488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_170
timestamp 1698175906
transform 1 0 20384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698175906
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_179
timestamp 1698175906
transform 1 0 21392 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_192
timestamp 1698175906
transform 1 0 22848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_196
timestamp 1698175906
transform 1 0 23296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_219
timestamp 1698175906
transform 1 0 25872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_226
timestamp 1698175906
transform 1 0 26656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_230
timestamp 1698175906
transform 1 0 27104 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_234
timestamp 1698175906
transform 1 0 27552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_236
timestamp 1698175906
transform 1 0 27776 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698175906
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_259
timestamp 1698175906
transform 1 0 30352 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_263
timestamp 1698175906
transform 1 0 30800 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_270
timestamp 1698175906
transform 1 0 31584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_274
timestamp 1698175906
transform 1 0 32032 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_306
timestamp 1698175906
transform 1 0 35616 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698175906
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_333
timestamp 1698175906
transform 1 0 38640 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_337
timestamp 1698175906
transform 1 0 39088 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_339
timestamp 1698175906
transform 1 0 39312 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_342
timestamp 1698175906
transform 1 0 39648 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_352
timestamp 1698175906
transform 1 0 40768 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_360
timestamp 1698175906
transform 1 0 41664 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_366
timestamp 1698175906
transform 1 0 42336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_370
timestamp 1698175906
transform 1 0 42784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698175906
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_394
timestamp 1698175906
transform 1 0 45472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_398
timestamp 1698175906
transform 1 0 45920 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_430
timestamp 1698175906
transform 1 0 49504 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_446
timestamp 1698175906
transform 1 0 51296 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698175906
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_457
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_34
timestamp 1698175906
transform 1 0 5152 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_38
timestamp 1698175906
transform 1 0 5600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_53
timestamp 1698175906
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_57
timestamp 1698175906
transform 1 0 7728 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698175906
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698175906
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_81
timestamp 1698175906
transform 1 0 10416 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_97
timestamp 1698175906
transform 1 0 12208 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_107
timestamp 1698175906
transform 1 0 13328 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_123
timestamp 1698175906
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698175906
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_192
timestamp 1698175906
transform 1 0 22848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_220
timestamp 1698175906
transform 1 0 25984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_224
timestamp 1698175906
transform 1 0 26432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_228
timestamp 1698175906
transform 1 0 26880 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_237
timestamp 1698175906
transform 1 0 27888 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_241
timestamp 1698175906
transform 1 0 28336 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_257
timestamp 1698175906
transform 1 0 30128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_270
timestamp 1698175906
transform 1 0 31584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_274
timestamp 1698175906
transform 1 0 32032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698175906
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_286
timestamp 1698175906
transform 1 0 33376 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_297
timestamp 1698175906
transform 1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_301
timestamp 1698175906
transform 1 0 35056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_305
timestamp 1698175906
transform 1 0 35504 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_337
timestamp 1698175906
transform 1 0 39088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698175906
transform 1 0 39984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698175906
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_368
timestamp 1698175906
transform 1 0 42560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_376
timestamp 1698175906
transform 1 0 43456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_378
timestamp 1698175906
transform 1 0 43680 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_381
timestamp 1698175906
transform 1 0 44016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_385
timestamp 1698175906
transform 1 0 44464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_395
timestamp 1698175906
transform 1 0 45584 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_411
timestamp 1698175906
transform 1 0 47376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698175906
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_430
timestamp 1698175906
transform 1 0 49504 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_18
timestamp 1698175906
transform 1 0 3360 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_26
timestamp 1698175906
transform 1 0 4256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_28
timestamp 1698175906
transform 1 0 4480 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_51
timestamp 1698175906
transform 1 0 7056 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_61
timestamp 1698175906
transform 1 0 8176 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_69
timestamp 1698175906
transform 1 0 9072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_71
timestamp 1698175906
transform 1 0 9296 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698175906
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_119
timestamp 1698175906
transform 1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_153
timestamp 1698175906
transform 1 0 18480 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_169
timestamp 1698175906
transform 1 0 20272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698175906
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_193
timestamp 1698175906
transform 1 0 22960 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_197
timestamp 1698175906
transform 1 0 23408 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_214
timestamp 1698175906
transform 1 0 25312 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_218
timestamp 1698175906
transform 1 0 25760 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_227
timestamp 1698175906
transform 1 0 26768 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_251
timestamp 1698175906
transform 1 0 29456 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_259
timestamp 1698175906
transform 1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_261
timestamp 1698175906
transform 1 0 30576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_274
timestamp 1698175906
transform 1 0 32032 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_278
timestamp 1698175906
transform 1 0 32480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_288
timestamp 1698175906
transform 1 0 33600 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_290
timestamp 1698175906
transform 1 0 33824 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_298
timestamp 1698175906
transform 1 0 34720 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698175906
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_321
timestamp 1698175906
transform 1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698175906
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_329
timestamp 1698175906
transform 1 0 38192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_338
timestamp 1698175906
transform 1 0 39200 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_373
timestamp 1698175906
transform 1 0 43120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_377
timestamp 1698175906
transform 1 0 43568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698175906
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_391
timestamp 1698175906
transform 1 0 45136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_393
timestamp 1698175906
transform 1 0 45360 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_423
timestamp 1698175906
transform 1 0 48720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_427
timestamp 1698175906
transform 1 0 49168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_431
timestamp 1698175906
transform 1 0 49616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_441
timestamp 1698175906
transform 1 0 50736 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_449
timestamp 1698175906
transform 1 0 51632 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_453
timestamp 1698175906
transform 1 0 52080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698175906
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_35
timestamp 1698175906
transform 1 0 5264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_68
timestamp 1698175906
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_76
timestamp 1698175906
transform 1 0 9856 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_108
timestamp 1698175906
transform 1 0 13440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_116
timestamp 1698175906
transform 1 0 14336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_118
timestamp 1698175906
transform 1 0 14560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_137
timestamp 1698175906
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698175906
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_174
timestamp 1698175906
transform 1 0 20832 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_178
timestamp 1698175906
transform 1 0 21280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_180
timestamp 1698175906
transform 1 0 21504 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_186
timestamp 1698175906
transform 1 0 22176 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_202
timestamp 1698175906
transform 1 0 23968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_227
timestamp 1698175906
transform 1 0 26768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_231
timestamp 1698175906
transform 1 0 27216 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_263
timestamp 1698175906
transform 1 0 30800 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698175906
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_284
timestamp 1698175906
transform 1 0 33152 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_330
timestamp 1698175906
transform 1 0 38304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698175906
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_352
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_369
timestamp 1698175906
transform 1 0 42672 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_373
timestamp 1698175906
transform 1 0 43120 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_387
timestamp 1698175906
transform 1 0 44688 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_393
timestamp 1698175906
transform 1 0 45360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_397
timestamp 1698175906
transform 1 0 45808 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_413
timestamp 1698175906
transform 1 0 47600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_417
timestamp 1698175906
transform 1 0 48048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698175906
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_433
timestamp 1698175906
transform 1 0 49840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_435
timestamp 1698175906
transform 1 0 50064 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_53
timestamp 1698175906
transform 1 0 7280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_57
timestamp 1698175906
transform 1 0 7728 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_64
timestamp 1698175906
transform 1 0 8512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_68
timestamp 1698175906
transform 1 0 8960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_90
timestamp 1698175906
transform 1 0 11424 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_98
timestamp 1698175906
transform 1 0 12320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_102
timestamp 1698175906
transform 1 0 12768 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_115
timestamp 1698175906
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_119
timestamp 1698175906
transform 1 0 14672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_146
timestamp 1698175906
transform 1 0 17696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_150
timestamp 1698175906
transform 1 0 18144 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_166
timestamp 1698175906
transform 1 0 19936 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698175906
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_181
timestamp 1698175906
transform 1 0 21616 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_190
timestamp 1698175906
transform 1 0 22624 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1698175906
transform 1 0 24416 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_208
timestamp 1698175906
transform 1 0 24640 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_238
timestamp 1698175906
transform 1 0 28000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698175906
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698175906
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_279
timestamp 1698175906
transform 1 0 32592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_283
timestamp 1698175906
transform 1 0 33040 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_287
timestamp 1698175906
transform 1 0 33488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_289
timestamp 1698175906
transform 1 0 33712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_292
timestamp 1698175906
transform 1 0 34048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_296
timestamp 1698175906
transform 1 0 34496 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698175906
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698175906
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_321
timestamp 1698175906
transform 1 0 37296 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_337
timestamp 1698175906
transform 1 0 39088 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_341
timestamp 1698175906
transform 1 0 39536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_345
timestamp 1698175906
transform 1 0 39984 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_353
timestamp 1698175906
transform 1 0 40880 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_357
timestamp 1698175906
transform 1 0 41328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_377
timestamp 1698175906
transform 1 0 43568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_401
timestamp 1698175906
transform 1 0 46256 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_417
timestamp 1698175906
transform 1 0 48048 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_421
timestamp 1698175906
transform 1 0 48496 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_434
timestamp 1698175906
transform 1 0 49952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_438
timestamp 1698175906
transform 1 0 50400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_440
timestamp 1698175906
transform 1 0 50624 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_447
timestamp 1698175906
transform 1 0 51408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698175906
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_57
timestamp 1698175906
transform 1 0 7728 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_65
timestamp 1698175906
transform 1 0 8624 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_80
timestamp 1698175906
transform 1 0 10304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_82
timestamp 1698175906
transform 1 0 10528 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_162
timestamp 1698175906
transform 1 0 19488 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_170
timestamp 1698175906
transform 1 0 20384 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_259
timestamp 1698175906
transform 1 0 30352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_263
timestamp 1698175906
transform 1 0 30800 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698175906
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_289
timestamp 1698175906
transform 1 0 33712 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_301
timestamp 1698175906
transform 1 0 35056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_305
timestamp 1698175906
transform 1 0 35504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_309
timestamp 1698175906
transform 1 0 35952 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_325
timestamp 1698175906
transform 1 0 37744 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_337
timestamp 1698175906
transform 1 0 39088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_339
timestamp 1698175906
transform 1 0 39312 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_342
timestamp 1698175906
transform 1 0 39648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_352
timestamp 1698175906
transform 1 0 40768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_386
timestamp 1698175906
transform 1 0 44576 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_418
timestamp 1698175906
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_422
timestamp 1698175906
transform 1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_426
timestamp 1698175906
transform 1 0 49056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_430
timestamp 1698175906
transform 1 0 49504 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_31
timestamp 1698175906
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_45
timestamp 1698175906
transform 1 0 6384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_84
timestamp 1698175906
transform 1 0 10752 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_88
timestamp 1698175906
transform 1 0 11200 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_90
timestamp 1698175906
transform 1 0 11424 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_93
timestamp 1698175906
transform 1 0 11760 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_97
timestamp 1698175906
transform 1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_115
timestamp 1698175906
transform 1 0 14224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_119
timestamp 1698175906
transform 1 0 14672 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_121
timestamp 1698175906
transform 1 0 14896 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_148
timestamp 1698175906
transform 1 0 17920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_170
timestamp 1698175906
transform 1 0 20384 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_174
timestamp 1698175906
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_209
timestamp 1698175906
transform 1 0 24752 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_219
timestamp 1698175906
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_223
timestamp 1698175906
transform 1 0 26320 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_239
timestamp 1698175906
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_243
timestamp 1698175906
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_251
timestamp 1698175906
transform 1 0 29456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698175906
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_259
timestamp 1698175906
transform 1 0 30352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_295
timestamp 1698175906
transform 1 0 34384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698175906
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698175906
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_351
timestamp 1698175906
transform 1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_355
timestamp 1698175906
transform 1 0 41104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_357
timestamp 1698175906
transform 1 0 41328 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_371
timestamp 1698175906
transform 1 0 42896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_377
timestamp 1698175906
transform 1 0 43568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698175906
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_434
timestamp 1698175906
transform 1 0 49952 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_438
timestamp 1698175906
transform 1 0 50400 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_447
timestamp 1698175906
transform 1 0 51408 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_457
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_18
timestamp 1698175906
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_26
timestamp 1698175906
transform 1 0 4256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_30
timestamp 1698175906
transform 1 0 4704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_56
timestamp 1698175906
transform 1 0 7616 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_64
timestamp 1698175906
transform 1 0 8512 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_68
timestamp 1698175906
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_79
timestamp 1698175906
transform 1 0 10192 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_111
timestamp 1698175906
transform 1 0 13776 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_115
timestamp 1698175906
transform 1 0 14224 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_119
timestamp 1698175906
transform 1 0 14672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_121
timestamp 1698175906
transform 1 0 14896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_134
timestamp 1698175906
transform 1 0 16352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698175906
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_167
timestamp 1698175906
transform 1 0 20048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_171
timestamp 1698175906
transform 1 0 20496 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_179
timestamp 1698175906
transform 1 0 21392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_181
timestamp 1698175906
transform 1 0 21616 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_194
timestamp 1698175906
transform 1 0 23072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_198
timestamp 1698175906
transform 1 0 23520 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_202
timestamp 1698175906
transform 1 0 23968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_224
timestamp 1698175906
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698175906
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_232
timestamp 1698175906
transform 1 0 27328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_240
timestamp 1698175906
transform 1 0 28224 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_244
timestamp 1698175906
transform 1 0 28672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_246
timestamp 1698175906
transform 1 0 28896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_249
timestamp 1698175906
transform 1 0 29232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_253
timestamp 1698175906
transform 1 0 29680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_286
timestamp 1698175906
transform 1 0 33376 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_295
timestamp 1698175906
transform 1 0 34384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_299
timestamp 1698175906
transform 1 0 34832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_301
timestamp 1698175906
transform 1 0 35056 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_333
timestamp 1698175906
transform 1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_337
timestamp 1698175906
transform 1 0 39088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_341
timestamp 1698175906
transform 1 0 39536 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_344
timestamp 1698175906
transform 1 0 39872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_374
timestamp 1698175906
transform 1 0 43232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_376
timestamp 1698175906
transform 1 0 43456 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_386
timestamp 1698175906
transform 1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_390
timestamp 1698175906
transform 1 0 45024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_394
timestamp 1698175906
transform 1 0 45472 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_398
timestamp 1698175906
transform 1 0 45920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_402
timestamp 1698175906
transform 1 0 46368 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_418
timestamp 1698175906
transform 1 0 48160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_422
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_428
timestamp 1698175906
transform 1 0 49280 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_432
timestamp 1698175906
transform 1 0 49728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_18
timestamp 1698175906
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_26
timestamp 1698175906
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_30
timestamp 1698175906
transform 1 0 4704 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698175906
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_44
timestamp 1698175906
transform 1 0 6272 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_60
timestamp 1698175906
transform 1 0 8064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_68
timestamp 1698175906
transform 1 0 8960 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_81
timestamp 1698175906
transform 1 0 10416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_85
timestamp 1698175906
transform 1 0 10864 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_127
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_130
timestamp 1698175906
transform 1 0 15904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_134
timestamp 1698175906
transform 1 0 16352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_169
timestamp 1698175906
transform 1 0 20272 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 20720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_179
timestamp 1698175906
transform 1 0 21392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_222
timestamp 1698175906
transform 1 0 26208 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_238
timestamp 1698175906
transform 1 0 28000 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_242
timestamp 1698175906
transform 1 0 28448 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698175906
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698175906
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_329
timestamp 1698175906
transform 1 0 38192 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_341
timestamp 1698175906
transform 1 0 39536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_354
timestamp 1698175906
transform 1 0 40992 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_362
timestamp 1698175906
transform 1 0 41888 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_368
timestamp 1698175906
transform 1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_372
timestamp 1698175906
transform 1 0 43008 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_376
timestamp 1698175906
transform 1 0 43456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_382
timestamp 1698175906
transform 1 0 44128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_384
timestamp 1698175906
transform 1 0 44352 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_392
timestamp 1698175906
transform 1 0 45248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_431
timestamp 1698175906
transform 1 0 49616 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_447
timestamp 1698175906
transform 1 0 51408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_457
timestamp 1698175906
transform 1 0 52528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_31
timestamp 1698175906
transform 1 0 4816 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_45
timestamp 1698175906
transform 1 0 6384 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_57
timestamp 1698175906
transform 1 0 7728 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_65
timestamp 1698175906
transform 1 0 8624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_67
timestamp 1698175906
transform 1 0 8848 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_101
timestamp 1698175906
transform 1 0 12656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_103
timestamp 1698175906
transform 1 0 12880 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_160
timestamp 1698175906
transform 1 0 19264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_176
timestamp 1698175906
transform 1 0 21056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_180
timestamp 1698175906
transform 1 0 21504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_188
timestamp 1698175906
transform 1 0 22400 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_194
timestamp 1698175906
transform 1 0 23072 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_223
timestamp 1698175906
transform 1 0 26320 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_251
timestamp 1698175906
transform 1 0 29456 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_255
timestamp 1698175906
transform 1 0 29904 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_271
timestamp 1698175906
transform 1 0 31696 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 32592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_314
timestamp 1698175906
transform 1 0 36512 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_324
timestamp 1698175906
transform 1 0 37632 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_340
timestamp 1698175906
transform 1 0 39424 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_352
timestamp 1698175906
transform 1 0 40768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_368
timestamp 1698175906
transform 1 0 42560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_399
timestamp 1698175906
transform 1 0 46032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_403
timestamp 1698175906
transform 1 0 46480 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_411
timestamp 1698175906
transform 1 0 47376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_415
timestamp 1698175906
transform 1 0 47824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_417
timestamp 1698175906
transform 1 0 48048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698175906
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_424
timestamp 1698175906
transform 1 0 48832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_433
timestamp 1698175906
transform 1 0 49840 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_437
timestamp 1698175906
transform 1 0 50288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_37
timestamp 1698175906
transform 1 0 5488 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_45
timestamp 1698175906
transform 1 0 6384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_52
timestamp 1698175906
transform 1 0 7168 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_84
timestamp 1698175906
transform 1 0 10752 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_100
timestamp 1698175906
transform 1 0 12544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698175906
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698175906
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_177
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_209
timestamp 1698175906
transform 1 0 24752 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_225
timestamp 1698175906
transform 1 0 26544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_229
timestamp 1698175906
transform 1 0 26992 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_257
timestamp 1698175906
transform 1 0 30128 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_273
timestamp 1698175906
transform 1 0 31920 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1698175906
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698175906
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_321
timestamp 1698175906
transform 1 0 37296 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_323
timestamp 1698175906
transform 1 0 37520 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_330
timestamp 1698175906
transform 1 0 38304 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_334
timestamp 1698175906
transform 1 0 38752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_336
timestamp 1698175906
transform 1 0 38976 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_366
timestamp 1698175906
transform 1 0 42336 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_370
timestamp 1698175906
transform 1 0 42784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_378
timestamp 1698175906
transform 1 0 43680 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_382
timestamp 1698175906
transform 1 0 44128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698175906
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_387
timestamp 1698175906
transform 1 0 44688 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_419
timestamp 1698175906
transform 1 0 48272 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_427
timestamp 1698175906
transform 1 0 49168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_431
timestamp 1698175906
transform 1 0 49616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_433
timestamp 1698175906
transform 1 0 49840 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_436
timestamp 1698175906
transform 1 0 50176 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_452
timestamp 1698175906
transform 1 0 51968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_454
timestamp 1698175906
transform 1 0 52192 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1698175906
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_34
timestamp 1698175906
transform 1 0 5152 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_42
timestamp 1698175906
transform 1 0 6048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_44
timestamp 1698175906
transform 1 0 6272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_53
timestamp 1698175906
transform 1 0 7280 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698175906
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_80
timestamp 1698175906
transform 1 0 10304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_84
timestamp 1698175906
transform 1 0 10752 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_92
timestamp 1698175906
transform 1 0 11648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_123
timestamp 1698175906
transform 1 0 15120 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_127
timestamp 1698175906
transform 1 0 15568 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_135
timestamp 1698175906
transform 1 0 16464 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698175906
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698175906
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_146
timestamp 1698175906
transform 1 0 17696 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_178
timestamp 1698175906
transform 1 0 21280 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_194
timestamp 1698175906
transform 1 0 23072 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_198
timestamp 1698175906
transform 1 0 23520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_200
timestamp 1698175906
transform 1 0 23744 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698175906
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_212
timestamp 1698175906
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_220
timestamp 1698175906
transform 1 0 25984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_224
timestamp 1698175906
transform 1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_226
timestamp 1698175906
transform 1 0 26656 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_239
timestamp 1698175906
transform 1 0 28112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_243
timestamp 1698175906
transform 1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_245
timestamp 1698175906
transform 1 0 28784 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_286
timestamp 1698175906
transform 1 0 33376 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_333
timestamp 1698175906
transform 1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_337
timestamp 1698175906
transform 1 0 39088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_360
timestamp 1698175906
transform 1 0 41664 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_376
timestamp 1698175906
transform 1 0 43456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_393
timestamp 1698175906
transform 1 0 45360 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_409
timestamp 1698175906
transform 1 0 47152 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_417
timestamp 1698175906
transform 1 0 48048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_419
timestamp 1698175906
transform 1 0 48272 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_422
timestamp 1698175906
transform 1 0 48608 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_426
timestamp 1698175906
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698175906
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_66
timestamp 1698175906
transform 1 0 8736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_70
timestamp 1698175906
transform 1 0 9184 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_74
timestamp 1698175906
transform 1 0 9632 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_90
timestamp 1698175906
transform 1 0 11424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_94
timestamp 1698175906
transform 1 0 11872 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_102
timestamp 1698175906
transform 1 0 12768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698175906
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_121
timestamp 1698175906
transform 1 0 14896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_123
timestamp 1698175906
transform 1 0 15120 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_155
timestamp 1698175906
transform 1 0 18704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_159
timestamp 1698175906
transform 1 0 19152 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_177
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_220
timestamp 1698175906
transform 1 0 25984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_224
timestamp 1698175906
transform 1 0 26432 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_232
timestamp 1698175906
transform 1 0 27328 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_251
timestamp 1698175906
transform 1 0 29456 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698175906
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_261
timestamp 1698175906
transform 1 0 30576 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_264
timestamp 1698175906
transform 1 0 30912 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_280
timestamp 1698175906
transform 1 0 32704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_284
timestamp 1698175906
transform 1 0 33152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_291
timestamp 1698175906
transform 1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_295
timestamp 1698175906
transform 1 0 34384 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698175906
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698175906
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_392
timestamp 1698175906
transform 1 0 45248 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_396
timestamp 1698175906
transform 1 0 45696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_398
timestamp 1698175906
transform 1 0 45920 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_430
timestamp 1698175906
transform 1 0 49504 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_444
timestamp 1698175906
transform 1 0 51072 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_452
timestamp 1698175906
transform 1 0 51968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698175906
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1698175906
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698175906
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_80
timestamp 1698175906
transform 1 0 10304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_86
timestamp 1698175906
transform 1 0 10976 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_102
timestamp 1698175906
transform 1 0 12768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_110
timestamp 1698175906
transform 1 0 13664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_114
timestamp 1698175906
transform 1 0 14112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_116
timestamp 1698175906
transform 1 0 14336 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_119
timestamp 1698175906
transform 1 0 14672 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_135
timestamp 1698175906
transform 1 0 16464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698175906
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_150
timestamp 1698175906
transform 1 0 18144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_154
timestamp 1698175906
transform 1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_156
timestamp 1698175906
transform 1 0 18816 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_161
timestamp 1698175906
transform 1 0 19376 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_165
timestamp 1698175906
transform 1 0 19824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_205
timestamp 1698175906
transform 1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698175906
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_212
timestamp 1698175906
transform 1 0 25088 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_244
timestamp 1698175906
transform 1 0 28672 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_252
timestamp 1698175906
transform 1 0 29568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_270
timestamp 1698175906
transform 1 0 31584 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698175906
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698175906
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_288
timestamp 1698175906
transform 1 0 33600 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_297
timestamp 1698175906
transform 1 0 34608 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_305
timestamp 1698175906
transform 1 0 35504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_336
timestamp 1698175906
transform 1 0 38976 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_340
timestamp 1698175906
transform 1 0 39424 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_348
timestamp 1698175906
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_358
timestamp 1698175906
transform 1 0 41440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_365
timestamp 1698175906
transform 1 0 42224 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_381
timestamp 1698175906
transform 1 0 44016 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_397
timestamp 1698175906
transform 1 0 45808 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_413
timestamp 1698175906
transform 1 0 47600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_417
timestamp 1698175906
transform 1 0 48048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698175906
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_422
timestamp 1698175906
transform 1 0 48608 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_438
timestamp 1698175906
transform 1 0 50400 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_45
timestamp 1698175906
transform 1 0 6384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_49
timestamp 1698175906
transform 1 0 6832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_51
timestamp 1698175906
transform 1 0 7056 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_81
timestamp 1698175906
transform 1 0 10416 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_89
timestamp 1698175906
transform 1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_93
timestamp 1698175906
transform 1 0 11760 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_97
timestamp 1698175906
transform 1 0 12208 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_117
timestamp 1698175906
transform 1 0 14448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_121
timestamp 1698175906
transform 1 0 14896 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_137
timestamp 1698175906
transform 1 0 16688 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_161
timestamp 1698175906
transform 1 0 19376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698175906
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_184
timestamp 1698175906
transform 1 0 21952 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_194
timestamp 1698175906
transform 1 0 23072 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_210
timestamp 1698175906
transform 1 0 24864 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_218
timestamp 1698175906
transform 1 0 25760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_222
timestamp 1698175906
transform 1 0 26208 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_238
timestamp 1698175906
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698175906
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698175906
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_247
timestamp 1698175906
transform 1 0 29008 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_255
timestamp 1698175906
transform 1 0 29904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_286
timestamp 1698175906
transform 1 0 33376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_296
timestamp 1698175906
transform 1 0 34496 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698175906
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698175906
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_330
timestamp 1698175906
transform 1 0 38304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_334
timestamp 1698175906
transform 1 0 38752 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_338
timestamp 1698175906
transform 1 0 39200 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_374
timestamp 1698175906
transform 1 0 43232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_378
timestamp 1698175906
transform 1 0 43680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_395
timestamp 1698175906
transform 1 0 45584 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_411
timestamp 1698175906
transform 1 0 47376 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_419
timestamp 1698175906
transform 1 0 48272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_457
timestamp 1698175906
transform 1 0 52528 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698175906
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_76
timestamp 1698175906
transform 1 0 9856 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_90
timestamp 1698175906
transform 1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_94
timestamp 1698175906
transform 1 0 11872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_110
timestamp 1698175906
transform 1 0 13664 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_126
timestamp 1698175906
transform 1 0 15456 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_134
timestamp 1698175906
transform 1 0 16352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698175906
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_174
timestamp 1698175906
transform 1 0 20832 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_182
timestamp 1698175906
transform 1 0 21728 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_186
timestamp 1698175906
transform 1 0 22176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698175906
transform 1 0 22624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_220
timestamp 1698175906
transform 1 0 25984 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_252
timestamp 1698175906
transform 1 0 29568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_256
timestamp 1698175906
transform 1 0 30016 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_272
timestamp 1698175906
transform 1 0 31808 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_284
timestamp 1698175906
transform 1 0 33152 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698175906
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_292
timestamp 1698175906
transform 1 0 34048 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_303
timestamp 1698175906
transform 1 0 35280 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_335
timestamp 1698175906
transform 1 0 38864 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_343
timestamp 1698175906
transform 1 0 39760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_347
timestamp 1698175906
transform 1 0 40208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698175906
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_352
timestamp 1698175906
transform 1 0 40768 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_361
timestamp 1698175906
transform 1 0 41776 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_377
timestamp 1698175906
transform 1 0 43568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_414
timestamp 1698175906
transform 1 0 47712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_418
timestamp 1698175906
transform 1 0 48160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_422
timestamp 1698175906
transform 1 0 48608 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_69
timestamp 1698175906
transform 1 0 9072 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_77
timestamp 1698175906
transform 1 0 9968 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_83
timestamp 1698175906
transform 1 0 10640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_87
timestamp 1698175906
transform 1 0 11088 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_95
timestamp 1698175906
transform 1 0 11984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_97
timestamp 1698175906
transform 1 0 12208 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698175906
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_107
timestamp 1698175906
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_115
timestamp 1698175906
transform 1 0 14224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_117
timestamp 1698175906
transform 1 0 14448 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_147
timestamp 1698175906
transform 1 0 17808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_151
timestamp 1698175906
transform 1 0 18256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_155
timestamp 1698175906
transform 1 0 18704 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_161
timestamp 1698175906
transform 1 0 19376 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_169
timestamp 1698175906
transform 1 0 20272 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_173
timestamp 1698175906
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_177
timestamp 1698175906
transform 1 0 21168 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_193
timestamp 1698175906
transform 1 0 22960 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_218
timestamp 1698175906
transform 1 0 25760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_228
timestamp 1698175906
transform 1 0 26880 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_232
timestamp 1698175906
transform 1 0 27328 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_235
timestamp 1698175906
transform 1 0 27664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_255
timestamp 1698175906
transform 1 0 29904 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_271
timestamp 1698175906
transform 1 0 31696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_275
timestamp 1698175906
transform 1 0 32144 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_278
timestamp 1698175906
transform 1 0 32480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_282
timestamp 1698175906
transform 1 0 32928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_286
timestamp 1698175906
transform 1 0 33376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_292
timestamp 1698175906
transform 1 0 34048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_296
timestamp 1698175906
transform 1 0 34496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_300
timestamp 1698175906
transform 1 0 34944 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_304
timestamp 1698175906
transform 1 0 35392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_306
timestamp 1698175906
transform 1 0 35616 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_312
timestamp 1698175906
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698175906
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_325
timestamp 1698175906
transform 1 0 37744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_327
timestamp 1698175906
transform 1 0 37968 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_334
timestamp 1698175906
transform 1 0 38752 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_347
timestamp 1698175906
transform 1 0 40208 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_379
timestamp 1698175906
transform 1 0 43792 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698175906
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_387
timestamp 1698175906
transform 1 0 44688 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_403
timestamp 1698175906
transform 1 0 46480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_436
timestamp 1698175906
transform 1 0 50176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_438
timestamp 1698175906
transform 1 0 50400 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_445
timestamp 1698175906
transform 1 0 51184 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_453
timestamp 1698175906
transform 1 0 52080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_457
timestamp 1698175906
transform 1 0 52528 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698175906
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_72
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_81
timestamp 1698175906
transform 1 0 10416 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_89
timestamp 1698175906
transform 1 0 11312 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_121
timestamp 1698175906
transform 1 0 14896 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_129
timestamp 1698175906
transform 1 0 15792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_131
timestamp 1698175906
transform 1 0 16016 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_146
timestamp 1698175906
transform 1 0 17696 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_154
timestamp 1698175906
transform 1 0 18592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_158
timestamp 1698175906
transform 1 0 19040 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_172
timestamp 1698175906
transform 1 0 20608 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_176
timestamp 1698175906
transform 1 0 21056 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_183
timestamp 1698175906
transform 1 0 21840 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_193
timestamp 1698175906
transform 1 0 22960 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698175906
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_212
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_244
timestamp 1698175906
transform 1 0 28672 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_247
timestamp 1698175906
transform 1 0 29008 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_263
timestamp 1698175906
transform 1 0 30800 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_267
timestamp 1698175906
transform 1 0 31248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698175906
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_290
timestamp 1698175906
transform 1 0 33824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698175906
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_354
timestamp 1698175906
transform 1 0 40992 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_365
timestamp 1698175906
transform 1 0 42224 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_381
timestamp 1698175906
transform 1 0 44016 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_387
timestamp 1698175906
transform 1 0 44688 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_403
timestamp 1698175906
transform 1 0 46480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_415
timestamp 1698175906
transform 1 0 47824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_419
timestamp 1698175906
transform 1 0 48272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_422
timestamp 1698175906
transform 1 0 48608 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_438
timestamp 1698175906
transform 1 0 50400 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_37
timestamp 1698175906
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_45
timestamp 1698175906
transform 1 0 6384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_76
timestamp 1698175906
transform 1 0 9856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_80
timestamp 1698175906
transform 1 0 10304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_121
timestamp 1698175906
transform 1 0 14896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_125
timestamp 1698175906
transform 1 0 15344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_127
timestamp 1698175906
transform 1 0 15568 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_136
timestamp 1698175906
transform 1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_140
timestamp 1698175906
transform 1 0 17024 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_149
timestamp 1698175906
transform 1 0 18032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_157
timestamp 1698175906
transform 1 0 18928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_169
timestamp 1698175906
transform 1 0 20272 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_173
timestamp 1698175906
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_214
timestamp 1698175906
transform 1 0 25312 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_224
timestamp 1698175906
transform 1 0 26432 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_240
timestamp 1698175906
transform 1 0 28224 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698175906
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_338
timestamp 1698175906
transform 1 0 39200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_353
timestamp 1698175906
transform 1 0 40880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_355
timestamp 1698175906
transform 1 0 41104 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_402
timestamp 1698175906
transform 1 0 46368 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_416
timestamp 1698175906
transform 1 0 47936 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_432
timestamp 1698175906
transform 1 0 49728 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698175906
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_457
timestamp 1698175906
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698175906
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_80
timestamp 1698175906
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_118
timestamp 1698175906
transform 1 0 14560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_122
timestamp 1698175906
transform 1 0 15008 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698175906
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_147
timestamp 1698175906
transform 1 0 17808 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_151
timestamp 1698175906
transform 1 0 18256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_153
timestamp 1698175906
transform 1 0 18480 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_170
timestamp 1698175906
transform 1 0 20384 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_198
timestamp 1698175906
transform 1 0 23520 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_206
timestamp 1698175906
transform 1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698175906
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_250
timestamp 1698175906
transform 1 0 29344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_254
timestamp 1698175906
transform 1 0 29792 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_262
timestamp 1698175906
transform 1 0 30688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_266
timestamp 1698175906
transform 1 0 31136 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_268
timestamp 1698175906
transform 1 0 31360 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_279
timestamp 1698175906
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_297
timestamp 1698175906
transform 1 0 34608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_327
timestamp 1698175906
transform 1 0 37968 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_337
timestamp 1698175906
transform 1 0 39088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_341
timestamp 1698175906
transform 1 0 39536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698175906
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698175906
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_359
timestamp 1698175906
transform 1 0 41552 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_361
timestamp 1698175906
transform 1 0 41776 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_370
timestamp 1698175906
transform 1 0 42784 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_406
timestamp 1698175906
transform 1 0 46816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_410
timestamp 1698175906
transform 1 0 47264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_426
timestamp 1698175906
transform 1 0 49056 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_69
timestamp 1698175906
transform 1 0 9072 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_77
timestamp 1698175906
transform 1 0 9968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_79
timestamp 1698175906
transform 1 0 10192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_88
timestamp 1698175906
transform 1 0 11200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_92
timestamp 1698175906
transform 1 0 11648 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_100
timestamp 1698175906
transform 1 0 12544 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698175906
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_123
timestamp 1698175906
transform 1 0 15120 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698175906
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_150
timestamp 1698175906
transform 1 0 18144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_154
timestamp 1698175906
transform 1 0 18592 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_170
timestamp 1698175906
transform 1 0 20384 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698175906
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698175906
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_179
timestamp 1698175906
transform 1 0 21392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_197
timestamp 1698175906
transform 1 0 23408 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_201
timestamp 1698175906
transform 1 0 23856 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_221
timestamp 1698175906
transform 1 0 26096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_225
timestamp 1698175906
transform 1 0 26544 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698175906
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_247
timestamp 1698175906
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_279
timestamp 1698175906
transform 1 0 32592 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_295
timestamp 1698175906
transform 1 0 34384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_303
timestamp 1698175906
transform 1 0 35280 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698175906
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_325
timestamp 1698175906
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_329
timestamp 1698175906
transform 1 0 38192 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_361
timestamp 1698175906
transform 1 0 41776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_374
timestamp 1698175906
transform 1 0 43232 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_382
timestamp 1698175906
transform 1 0 44128 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_435
timestamp 1698175906
transform 1 0 50064 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698175906
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_457
timestamp 1698175906
transform 1 0 52528 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698175906
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_72
timestamp 1698175906
transform 1 0 9408 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_88
timestamp 1698175906
transform 1 0 11200 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_96
timestamp 1698175906
transform 1 0 12096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_100
timestamp 1698175906
transform 1 0 12544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698175906
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_146
timestamp 1698175906
transform 1 0 17696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_150
timestamp 1698175906
transform 1 0 18144 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_158
timestamp 1698175906
transform 1 0 19040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_162
timestamp 1698175906
transform 1 0 19488 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_166
timestamp 1698175906
transform 1 0 19936 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_168
timestamp 1698175906
transform 1 0 20160 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_178
timestamp 1698175906
transform 1 0 21280 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_186
timestamp 1698175906
transform 1 0 22176 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_190
timestamp 1698175906
transform 1 0 22624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_192
timestamp 1698175906
transform 1 0 22848 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_201
timestamp 1698175906
transform 1 0 23856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_205
timestamp 1698175906
transform 1 0 24304 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698175906
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_212
timestamp 1698175906
transform 1 0 25088 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_220
timestamp 1698175906
transform 1 0 25984 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_229
timestamp 1698175906
transform 1 0 26992 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_233
timestamp 1698175906
transform 1 0 27440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_235
timestamp 1698175906
transform 1 0 27664 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_265
timestamp 1698175906
transform 1 0 31024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_269
timestamp 1698175906
transform 1 0 31472 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_273
timestamp 1698175906
transform 1 0 31920 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_277
timestamp 1698175906
transform 1 0 32368 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698175906
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_288
timestamp 1698175906
transform 1 0 33600 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_304
timestamp 1698175906
transform 1 0 35392 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_308
timestamp 1698175906
transform 1 0 35840 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_310
timestamp 1698175906
transform 1 0 36064 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_352
timestamp 1698175906
transform 1 0 40768 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_367
timestamp 1698175906
transform 1 0 42448 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_403
timestamp 1698175906
transform 1 0 46480 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_411
timestamp 1698175906
transform 1 0 47376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_418
timestamp 1698175906
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_422
timestamp 1698175906
transform 1 0 48608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_430
timestamp 1698175906
transform 1 0 49504 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_434
timestamp 1698175906
transform 1 0 49952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_69
timestamp 1698175906
transform 1 0 9072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_102
timestamp 1698175906
transform 1 0 12768 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1698175906
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_107
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_123
timestamp 1698175906
transform 1 0 15120 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_166
timestamp 1698175906
transform 1 0 19936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_185
timestamp 1698175906
transform 1 0 22064 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_201
timestamp 1698175906
transform 1 0 23856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_211
timestamp 1698175906
transform 1 0 24976 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_215
timestamp 1698175906
transform 1 0 25424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_217
timestamp 1698175906
transform 1 0 25648 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_224
timestamp 1698175906
transform 1 0 26432 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_232
timestamp 1698175906
transform 1 0 27328 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_242
timestamp 1698175906
transform 1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698175906
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_247
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_263
timestamp 1698175906
transform 1 0 30800 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_300
timestamp 1698175906
transform 1 0 34944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_304
timestamp 1698175906
transform 1 0 35392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_312
timestamp 1698175906
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698175906
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_328
timestamp 1698175906
transform 1 0 38080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_332
timestamp 1698175906
transform 1 0 38528 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_342
timestamp 1698175906
transform 1 0 39648 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_358
timestamp 1698175906
transform 1 0 41440 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_362
timestamp 1698175906
transform 1 0 41888 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_364
timestamp 1698175906
transform 1 0 42112 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_374
timestamp 1698175906
transform 1 0 43232 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_382
timestamp 1698175906
transform 1 0 44128 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_384
timestamp 1698175906
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_387
timestamp 1698175906
transform 1 0 44688 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_403
timestamp 1698175906
transform 1 0 46480 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_405
timestamp 1698175906
transform 1 0 46704 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_408
timestamp 1698175906
transform 1 0 47040 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_416
timestamp 1698175906
transform 1 0 47936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_420
timestamp 1698175906
transform 1 0 48384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_446
timestamp 1698175906
transform 1 0 51296 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698175906
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_457
timestamp 1698175906
transform 1 0 52528 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698175906
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698175906
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698175906
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698175906
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_212
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_216
timestamp 1698175906
transform 1 0 25536 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_221
timestamp 1698175906
transform 1 0 26096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_225
timestamp 1698175906
transform 1 0 26544 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_257
timestamp 1698175906
transform 1 0 30128 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_273
timestamp 1698175906
transform 1 0 31920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698175906
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698175906
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_282
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_290
timestamp 1698175906
transform 1 0 33824 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_303
timestamp 1698175906
transform 1 0 35280 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_341
timestamp 1698175906
transform 1 0 39536 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698175906
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_352
timestamp 1698175906
transform 1 0 40768 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_384
timestamp 1698175906
transform 1 0 44352 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_392
timestamp 1698175906
transform 1 0 45248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_396
timestamp 1698175906
transform 1 0 45696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_416
timestamp 1698175906
transform 1 0 47936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_432
timestamp 1698175906
transform 1 0 49728 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_436
timestamp 1698175906
transform 1 0 50176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_438
timestamp 1698175906
transform 1 0 50400 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698175906
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_139
timestamp 1698175906
transform 1 0 16912 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_155
timestamp 1698175906
transform 1 0 18704 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_163
timestamp 1698175906
transform 1 0 19600 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_167
timestamp 1698175906
transform 1 0 20048 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_204
timestamp 1698175906
transform 1 0 24192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_208
timestamp 1698175906
transform 1 0 24640 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_227
timestamp 1698175906
transform 1 0 26768 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_231
timestamp 1698175906
transform 1 0 27216 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_239
timestamp 1698175906
transform 1 0 28112 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_243
timestamp 1698175906
transform 1 0 28560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698175906
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698175906
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_349
timestamp 1698175906
transform 1 0 40432 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_357
timestamp 1698175906
transform 1 0 41328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_361
timestamp 1698175906
transform 1 0 41776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_363
timestamp 1698175906
transform 1 0 42000 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_372
timestamp 1698175906
transform 1 0 43008 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_380
timestamp 1698175906
transform 1 0 43904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698175906
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_387
timestamp 1698175906
transform 1 0 44688 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_395
timestamp 1698175906
transform 1 0 45584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_406
timestamp 1698175906
transform 1 0 46816 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_414
timestamp 1698175906
transform 1 0 47712 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_418
timestamp 1698175906
transform 1 0 48160 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_457
timestamp 1698175906
transform 1 0 52528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698175906
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698175906
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698175906
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698175906
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_142
timestamp 1698175906
transform 1 0 17248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_158
timestamp 1698175906
transform 1 0 19040 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_172
timestamp 1698175906
transform 1 0 20608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_174
timestamp 1698175906
transform 1 0 20832 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_180
timestamp 1698175906
transform 1 0 21504 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_187
timestamp 1698175906
transform 1 0 22288 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_191
timestamp 1698175906
transform 1 0 22736 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_193
timestamp 1698175906
transform 1 0 22960 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_200
timestamp 1698175906
transform 1 0 23744 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698175906
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_212
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_216
timestamp 1698175906
transform 1 0 25536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_236
timestamp 1698175906
transform 1 0 27776 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_240
timestamp 1698175906
transform 1 0 28224 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698175906
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698175906
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_282
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_286
timestamp 1698175906
transform 1 0 33376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_303
timestamp 1698175906
transform 1 0 35280 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_311
timestamp 1698175906
transform 1 0 36176 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_328
timestamp 1698175906
transform 1 0 38080 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_336
timestamp 1698175906
transform 1 0 38976 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698175906
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_358
timestamp 1698175906
transform 1 0 41440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_397
timestamp 1698175906
transform 1 0 45808 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_413
timestamp 1698175906
transform 1 0 47600 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1698175906
transform 1 0 48048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698175906
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_422
timestamp 1698175906
transform 1 0 48608 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698175906
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698175906
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698175906
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698175906
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_123
timestamp 1698175906
transform 1 0 15120 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_131
timestamp 1698175906
transform 1 0 16016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_135
timestamp 1698175906
transform 1 0 16464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_166
timestamp 1698175906
transform 1 0 19936 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_170
timestamp 1698175906
transform 1 0 20384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698175906
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_185
timestamp 1698175906
transform 1 0 22064 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_189
timestamp 1698175906
transform 1 0 22512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_207
timestamp 1698175906
transform 1 0 24528 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_215
timestamp 1698175906
transform 1 0 25424 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_219
timestamp 1698175906
transform 1 0 25872 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_229
timestamp 1698175906
transform 1 0 26992 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_305
timestamp 1698175906
transform 1 0 35504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_309
timestamp 1698175906
transform 1 0 35952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698175906
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_375
timestamp 1698175906
transform 1 0 43344 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_383
timestamp 1698175906
transform 1 0 44240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_387
timestamp 1698175906
transform 1 0 44688 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_424
timestamp 1698175906
transform 1 0 48832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_428
timestamp 1698175906
transform 1 0 49280 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_457
timestamp 1698175906
transform 1 0 52528 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_2
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_36
timestamp 1698175906
transform 1 0 5376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_70
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_104
timestamp 1698175906
transform 1 0 12992 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_138
timestamp 1698175906
transform 1 0 16800 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_172
timestamp 1698175906
transform 1 0 20608 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_206
timestamp 1698175906
transform 1 0 24416 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_240
timestamp 1698175906
transform 1 0 28224 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_274
timestamp 1698175906
transform 1 0 32032 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_278
timestamp 1698175906
transform 1 0 32480 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_294
timestamp 1698175906
transform 1 0 34272 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_302
timestamp 1698175906
transform 1 0 35168 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_308
timestamp 1698175906
transform 1 0 35840 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_342
timestamp 1698175906
transform 1 0 39648 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_350
timestamp 1698175906
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_354
timestamp 1698175906
transform 1 0 40992 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_365
timestamp 1698175906
transform 1 0 42224 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_373
timestamp 1698175906
transform 1 0 43120 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_376
timestamp 1698175906
transform 1 0 43456 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_410
timestamp 1698175906
transform 1 0 47264 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_452
timestamp 1698175906
transform 1 0 51968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_460
timestamp 1698175906
transform 1 0 52864 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_464
timestamp 1698175906
transform 1 0 53312 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698175906
transform -1 0 53424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698175906
transform -1 0 53424 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698175906
transform -1 0 53424 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698175906
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698175906
transform -1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform -1 0 53424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698175906
transform -1 0 53424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform -1 0 53424 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698175906
transform -1 0 53424 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698175906
transform -1 0 53424 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform -1 0 53424 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698175906
transform -1 0 53424 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698175906
transform -1 0 53424 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 2800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input16
timestamp 1698175906
transform 1 0 41328 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 50512 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 50512 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 50512 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 49392 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 50512 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 50512 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 49392 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform -1 0 52304 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform -1 0 12096 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698175906
transform -1 0 14672 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698175906
transform -1 0 50848 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_62 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 53648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_63
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 53648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_64
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 53648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_65
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 53648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_66
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 53648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_67
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 53648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_68
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 53648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 53648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 53648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_72
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 53648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_73
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 53648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_74
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 53648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_75
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 53648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_76
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 53648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_77
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 53648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_78
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 53648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_79
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 53648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_80
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 53648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_81
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 53648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_82
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 53648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_83
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 53648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_84
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 53648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_85
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 53648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_86
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 53648 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_87
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 53648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_88
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 53648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_89
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 53648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_90
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 53648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_91
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 53648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_92
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 53648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_93
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 53648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_94
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 53648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_95
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 53648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_96
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 53648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_97
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 53648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_98
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 53648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_99
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 53648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_100
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 53648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_101
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 53648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_102
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 53648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_103
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 53648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_104
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 53648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_105
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 53648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_106
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 53648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_107
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 53648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_108
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 53648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_109
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 53648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_110
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 53648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_111
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 53648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_112
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 53648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_113
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 53648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_114
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 53648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_115
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 53648 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_116
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 53648 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_117
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 53648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_118
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 53648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_119
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 53648 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_120
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 53648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_121
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 53648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_122
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 53648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_123
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 53648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_30
timestamp 1698175906
transform -1 0 25648 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_31
timestamp 1698175906
transform -1 0 17248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  serial_ports_32 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_124 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_125
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_126
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_127
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_128
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_129
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_130
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_131
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_132
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_133
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_134
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_135
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_137
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_138
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_139
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_140
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_141
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_142
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_143
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_144
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_145
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_146
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_147
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_148
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_149
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_150
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_151
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_152
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_153
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_154
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_156
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_157
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_161
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_162
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_164
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_165
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_166
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_167
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_168
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_169
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_170
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_171
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_172
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_173
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_174
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_175
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_176
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_177
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_178
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_179
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_180
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_181
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_182
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_183
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_184
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_185
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_186
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_187
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_188
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_189
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_190
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_191
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_192
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_193
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_194
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_195
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_196
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_197
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_198
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_199
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_200
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_201
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_202
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_203
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_204
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_205
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_206
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_207
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_208
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_209
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_210
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_211
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_212
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_213
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_214
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_215
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_216
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_217
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_218
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_219
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_220
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_221
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_222
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_223
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_224
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_225
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_226
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_227
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_228
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_229
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_230
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_231
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_232
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_233
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_234
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_235
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_236
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_237
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_238
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_239
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_240
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_241
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_242
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_243
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_244
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_245
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_246
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_247
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_248
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_249
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_250
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_251
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_252
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_253
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_254
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_255
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_256
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_257
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_258
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_259
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_260
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_261
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_262
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_263
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_264
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_265
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_266
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_267
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_268
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_269
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_270
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_271
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_272
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_273
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_274
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_275
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_276
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_277
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_278
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_279
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_280
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_281
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_282
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_283
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_284
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_285
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_286
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_287
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_288
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_289
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_290
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_291
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_292
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_293
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_294
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_295
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_296
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_297
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_298
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_299
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_300
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_301
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_302
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_303
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_304
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_305
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_306
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_307
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_308
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_309
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_310
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_311
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_312
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_313
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_314
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_315
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_316
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_317
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_318
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_319
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_320
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_321
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_322
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_323
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_324
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_325
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_326
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_327
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_328
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_329
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_330
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_331
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_332
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_333
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_334
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_335
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_336
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_337
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_338
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_339
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_340
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_341
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_342
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_343
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_344
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_345
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_346
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_347
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_348
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_349
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_350
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_351
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_352
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_353
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_354
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_355
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_356
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_357
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_358
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_359
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_360
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_361
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_362
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_363
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_364
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_365
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_366
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_367
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_368
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_369
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_370
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_371
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_372
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_373
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_374
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_375
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_376
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_377
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_378
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_379
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_380
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_381
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_382
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_383
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_384
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_385
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_386
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_387
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_388
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_389
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_390
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_391
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_392
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_393
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_394
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_395
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_396
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_397
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_398
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_399
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_400
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_401
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_402
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_403
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_404
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_405
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_406
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_407
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_408
timestamp 1698175906
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_409
timestamp 1698175906
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_410
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_411
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_412
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_413
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_414
timestamp 1698175906
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_415
timestamp 1698175906
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_416
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_417
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_418
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_419
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_420
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_421
timestamp 1698175906
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_422
timestamp 1698175906
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_423
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_424
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_425
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_426
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_427
timestamp 1698175906
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_428
timestamp 1698175906
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_429
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_430
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_431
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_432
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_433
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_434
timestamp 1698175906
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_435
timestamp 1698175906
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_436
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_437
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_438
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_439
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_440
timestamp 1698175906
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_441
timestamp 1698175906
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_442
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_443
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_444
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_445
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_446
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_447
timestamp 1698175906
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_448
timestamp 1698175906
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_449
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_450
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_451
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_452
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_453
timestamp 1698175906
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_454
timestamp 1698175906
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_455
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_456
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_457
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_458
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_459
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_460
timestamp 1698175906
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_461
timestamp 1698175906
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_462
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_463
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_464
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_465
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_466
timestamp 1698175906
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_467
timestamp 1698175906
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_468
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_469
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_470
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_471
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_472
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_473
timestamp 1698175906
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_474
timestamp 1698175906
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_475
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_476
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_477
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_478
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_479
timestamp 1698175906
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_480
timestamp 1698175906
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_481
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_482
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_483
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_484
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_485
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_486
timestamp 1698175906
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_487
timestamp 1698175906
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_488
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_489
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_490
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_491
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_492
timestamp 1698175906
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_493
timestamp 1698175906
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_494
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_495
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_496
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_497
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_498
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_499
timestamp 1698175906
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_500
timestamp 1698175906
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_501
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_502
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_503
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_504
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_505
timestamp 1698175906
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_506
timestamp 1698175906
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_507
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_508
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_509
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_510
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_511
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_512
timestamp 1698175906
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_513
timestamp 1698175906
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_514
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_515
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_516
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_517
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_518
timestamp 1698175906
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_519
timestamp 1698175906
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_520
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_521
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_522
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_523
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_524
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_525
timestamp 1698175906
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_526
timestamp 1698175906
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_527
timestamp 1698175906
transform 1 0 5152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_528
timestamp 1698175906
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_529
timestamp 1698175906
transform 1 0 12768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_530
timestamp 1698175906
transform 1 0 16576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_531
timestamp 1698175906
transform 1 0 20384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_532
timestamp 1698175906
transform 1 0 24192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_533
timestamp 1698175906
transform 1 0 28000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_534
timestamp 1698175906
transform 1 0 31808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_535
timestamp 1698175906
transform 1 0 35616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_536
timestamp 1698175906
transform 1 0 39424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_537
timestamp 1698175906
transform 1 0 43232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_538
timestamp 1698175906
transform 1 0 47040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_539
timestamp 1698175906
transform 1 0 50848 0 -1 51744
box -86 -86 310 870
<< labels >>
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 RXD
port 0 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 TXD
port 1 nsew signal tristate
flabel metal3 s 54200 3136 55000 3248 0 FreeSans 448 0 0 0 addr[0]
port 2 nsew signal input
flabel metal3 s 54200 5824 55000 5936 0 FreeSans 448 0 0 0 addr[1]
port 3 nsew signal input
flabel metal3 s 54200 8512 55000 8624 0 FreeSans 448 0 0 0 addr[2]
port 4 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 bus_cyc
port 5 nsew signal input
flabel metal2 s 47488 0 47600 800 0 FreeSans 448 90 0 0 bus_we
port 6 nsew signal input
flabel metal3 s 54200 11200 55000 11312 0 FreeSans 448 0 0 0 data_in[0]
port 7 nsew signal input
flabel metal3 s 54200 13888 55000 14000 0 FreeSans 448 0 0 0 data_in[1]
port 8 nsew signal input
flabel metal3 s 54200 16576 55000 16688 0 FreeSans 448 0 0 0 data_in[2]
port 9 nsew signal input
flabel metal3 s 54200 19264 55000 19376 0 FreeSans 448 0 0 0 data_in[3]
port 10 nsew signal input
flabel metal3 s 54200 21952 55000 22064 0 FreeSans 448 0 0 0 data_in[4]
port 11 nsew signal input
flabel metal3 s 54200 24640 55000 24752 0 FreeSans 448 0 0 0 data_in[5]
port 12 nsew signal input
flabel metal3 s 54200 27328 55000 27440 0 FreeSans 448 0 0 0 data_in[6]
port 13 nsew signal input
flabel metal3 s 54200 30016 55000 30128 0 FreeSans 448 0 0 0 data_in[7]
port 14 nsew signal input
flabel metal3 s 54200 32704 55000 32816 0 FreeSans 448 0 0 0 data_out[0]
port 15 nsew signal tristate
flabel metal3 s 54200 35392 55000 35504 0 FreeSans 448 0 0 0 data_out[1]
port 16 nsew signal tristate
flabel metal3 s 54200 38080 55000 38192 0 FreeSans 448 0 0 0 data_out[2]
port 17 nsew signal tristate
flabel metal3 s 54200 40768 55000 40880 0 FreeSans 448 0 0 0 data_out[3]
port 18 nsew signal tristate
flabel metal3 s 54200 43456 55000 43568 0 FreeSans 448 0 0 0 data_out[4]
port 19 nsew signal tristate
flabel metal3 s 54200 46144 55000 46256 0 FreeSans 448 0 0 0 data_out[5]
port 20 nsew signal tristate
flabel metal3 s 54200 48832 55000 48944 0 FreeSans 448 0 0 0 data_out[6]
port 21 nsew signal tristate
flabel metal3 s 54200 51520 55000 51632 0 FreeSans 448 0 0 0 data_out[7]
port 22 nsew signal tristate
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_in
port 23 nsew signal input
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 24 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 25 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 26 nsew signal tristate
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 io_out[0]
port 27 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 io_out[1]
port 28 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 io_out[2]
port 29 nsew signal tristate
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 irq3
port 30 nsew signal tristate
flabel metal2 s 41216 54200 41328 55000 0 FreeSans 448 90 0 0 rst
port 31 nsew signal input
flabel metal4 s 4448 3076 4768 51804 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 35168 3076 35488 51804 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 19808 3076 20128 51804 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 51804 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal2 s 13664 54200 13776 55000 0 FreeSans 448 90 0 0 wb_clk_i
port 34 nsew signal input
rlabel metal1 27496 50960 27496 50960 0 vdd
rlabel metal1 27496 51744 27496 51744 0 vss
rlabel metal3 39592 3416 39592 3416 0 RXD
rlabel metal3 35560 3640 35560 3640 0 TXD
rlabel metal2 45360 20552 45360 20552 0 _0000_
rlabel metal2 46704 17752 46704 17752 0 _0001_
rlabel metal2 48888 14896 48888 14896 0 _0002_
rlabel metal2 51128 12880 51128 12880 0 _0003_
rlabel metal2 51072 18648 51072 18648 0 _0004_
rlabel metal2 52808 22736 52808 22736 0 _0005_
rlabel metal3 52080 27272 52080 27272 0 _0006_
rlabel metal2 46648 24360 46648 24360 0 _0007_
rlabel metal2 51128 10920 51128 10920 0 _0008_
rlabel metal2 51128 6216 51128 6216 0 _0009_
rlabel metal2 47488 4536 47488 4536 0 _0010_
rlabel metal2 44408 3864 44408 3864 0 _0011_
rlabel metal2 46984 11312 46984 11312 0 _0012_
rlabel metal2 26264 18760 26264 18760 0 _0013_
rlabel metal2 31640 8792 31640 8792 0 _0014_
rlabel metal2 31864 12600 31864 12600 0 _0015_
rlabel metal2 30576 14280 30576 14280 0 _0016_
rlabel metal3 43008 15176 43008 15176 0 _0017_
rlabel metal2 42616 13384 42616 13384 0 _0018_
rlabel metal2 34832 5992 34832 5992 0 _0019_
rlabel metal2 36232 5096 36232 5096 0 _0020_
rlabel metal2 38808 6440 38808 6440 0 _0021_
rlabel metal2 41944 5432 41944 5432 0 _0022_
rlabel metal2 27608 10920 27608 10920 0 _0023_
rlabel metal3 26768 13608 26768 13608 0 _0024_
rlabel metal2 23912 12992 23912 12992 0 _0025_
rlabel metal2 25704 15848 25704 15848 0 _0026_
rlabel metal2 23352 16296 23352 16296 0 _0027_
rlabel metal2 23576 21000 23576 21000 0 _0028_
rlabel metal2 23912 19600 23912 19600 0 _0029_
rlabel metal3 26320 22232 26320 22232 0 _0030_
rlabel metal2 31976 4760 31976 4760 0 _0031_
rlabel metal3 31864 25592 31864 25592 0 _0032_
rlabel metal3 29848 26936 29848 26936 0 _0033_
rlabel metal2 31080 32592 31080 32592 0 _0034_
rlabel metal2 32144 28728 32144 28728 0 _0035_
rlabel metal2 34720 31752 34720 31752 0 _0036_
rlabel metal2 33880 36512 33880 36512 0 _0037_
rlabel metal2 36120 38668 36120 38668 0 _0038_
rlabel metal2 35112 35224 35112 35224 0 _0039_
rlabel metal3 50568 4424 50568 4424 0 _0040_
rlabel metal2 52472 31472 52472 31472 0 _0041_
rlabel metal3 45976 35000 45976 35000 0 _0042_
rlabel metal3 46536 36568 46536 36568 0 _0043_
rlabel metal2 52472 32872 52472 32872 0 _0044_
rlabel metal2 51128 35280 51128 35280 0 _0045_
rlabel metal2 51072 42056 51072 42056 0 _0046_
rlabel metal2 51128 39312 51128 39312 0 _0047_
rlabel metal2 51800 44688 51800 44688 0 _0048_
rlabel metal2 46592 48440 46592 48440 0 _0049_
rlabel metal2 51128 47152 51128 47152 0 _0050_
rlabel metal2 51240 49896 51240 49896 0 _0051_
rlabel metal2 47824 42840 47824 42840 0 _0052_
rlabel metal3 49728 29512 49728 29512 0 _0053_
rlabel metal2 26264 24304 26264 24304 0 _0054_
rlabel metal2 29960 24528 29960 24528 0 _0055_
rlabel metal2 27272 32760 27272 32760 0 _0056_
rlabel metal2 26264 32984 26264 32984 0 _0057_
rlabel metal3 21056 31080 21056 31080 0 _0058_
rlabel metal2 22008 33488 22008 33488 0 _0059_
rlabel metal2 21560 26264 21560 26264 0 _0060_
rlabel metal3 23576 27160 23576 27160 0 _0061_
rlabel metal2 32648 23520 32648 23520 0 _0062_
rlabel metal2 36232 24304 36232 24304 0 _0063_
rlabel metal2 33656 18032 33656 18032 0 _0064_
rlabel metal2 29960 18032 29960 18032 0 _0065_
rlabel metal2 41160 30632 41160 30632 0 _0066_
rlabel metal2 37408 28616 37408 28616 0 _0067_
rlabel metal3 41496 26152 41496 26152 0 _0068_
rlabel metal3 41328 29288 41328 29288 0 _0069_
rlabel metal2 27048 42448 27048 42448 0 _0070_
rlabel metal2 18984 39144 18984 39144 0 _0071_
rlabel metal2 22792 40320 22792 40320 0 _0072_
rlabel metal2 16184 40320 16184 40320 0 _0073_
rlabel metal3 19544 50456 19544 50456 0 _0074_
rlabel metal3 29064 46760 29064 46760 0 _0075_
rlabel metal3 28840 50680 28840 50680 0 _0076_
rlabel metal3 29008 49672 29008 49672 0 _0077_
rlabel metal2 26320 44520 26320 44520 0 _0078_
rlabel metal3 19208 47320 19208 47320 0 _0079_
rlabel metal2 15512 43064 15512 43064 0 _0080_
rlabel metal3 15008 46536 15008 46536 0 _0081_
rlabel metal2 7560 43904 7560 43904 0 _0082_
rlabel metal2 10920 46648 10920 46648 0 _0083_
rlabel metal2 8120 41552 8120 41552 0 _0084_
rlabel metal3 13384 38920 13384 38920 0 _0085_
rlabel metal2 33096 46928 33096 46928 0 _0086_
rlabel metal3 33600 50456 33600 50456 0 _0087_
rlabel metal3 38416 50456 38416 50456 0 _0088_
rlabel metal2 41048 50232 41048 50232 0 _0089_
rlabel metal2 42280 49840 42280 49840 0 _0090_
rlabel metal3 43624 46536 43624 46536 0 _0091_
rlabel metal2 42280 44408 42280 44408 0 _0092_
rlabel metal2 37464 45584 37464 45584 0 _0093_
rlabel metal2 29792 42504 29792 42504 0 _0094_
rlabel metal2 2296 13216 2296 13216 0 _0095_
rlabel metal2 2520 11760 2520 11760 0 _0096_
rlabel metal2 2520 17024 2520 17024 0 _0097_
rlabel metal2 4312 10192 4312 10192 0 _0098_
rlabel metal2 6104 8232 6104 8232 0 _0099_
rlabel metal2 8120 8960 8120 8960 0 _0100_
rlabel metal2 11088 7560 11088 7560 0 _0101_
rlabel metal2 14280 7532 14280 7532 0 _0102_
rlabel metal2 15456 8344 15456 8344 0 _0103_
rlabel metal2 17416 10976 17416 10976 0 _0104_
rlabel metal2 19544 15456 19544 15456 0 _0105_
rlabel metal2 18648 17304 18648 17304 0 _0106_
rlabel metal2 13272 17696 13272 17696 0 _0107_
rlabel metal2 10416 15960 10416 15960 0 _0108_
rlabel metal3 13608 29288 13608 29288 0 _0109_
rlabel metal2 10136 31416 10136 31416 0 _0110_
rlabel metal3 13608 26936 13608 26936 0 _0111_
rlabel metal2 14728 24472 14728 24472 0 _0112_
rlabel metal2 6552 34552 6552 34552 0 _0113_
rlabel metal2 10024 36848 10024 36848 0 _0114_
rlabel metal3 4144 37128 4144 37128 0 _0115_
rlabel metal2 6888 39256 6888 39256 0 _0116_
rlabel metal2 2632 24360 2632 24360 0 _0117_
rlabel metal3 4704 27720 4704 27720 0 _0118_
rlabel metal3 4424 30072 4424 30072 0 _0119_
rlabel metal2 2520 32144 2520 32144 0 _0120_
rlabel metal2 2520 19544 2520 19544 0 _0121_
rlabel metal2 2632 21840 2632 21840 0 _0122_
rlabel metal2 10808 21504 10808 21504 0 _0123_
rlabel metal2 14280 21728 14280 21728 0 _0124_
rlabel metal2 45304 31416 45304 31416 0 _0125_
rlabel metal2 9688 6160 9688 6160 0 _0126_
rlabel metal2 28728 7784 28728 7784 0 _0127_
rlabel metal2 20720 10696 20720 10696 0 _0128_
rlabel metal2 20496 7560 20496 7560 0 _0129_
rlabel metal2 17752 6944 17752 6944 0 _0130_
rlabel metal2 19208 5152 19208 5152 0 _0131_
rlabel metal2 20776 4816 20776 4816 0 _0132_
rlabel metal2 25424 3640 25424 3640 0 _0133_
rlabel metal2 29960 4648 29960 4648 0 _0134_
rlabel metal2 9744 5208 9744 5208 0 _0135_
rlabel metal2 36680 40712 36680 40712 0 _0136_
rlabel metal2 30464 38920 30464 38920 0 _0137_
rlabel metal3 32480 41048 32480 41048 0 _0138_
rlabel metal2 40936 41328 40936 41328 0 _0139_
rlabel metal2 45080 41384 45080 41384 0 _0140_
rlabel metal2 48552 39984 48552 39984 0 _0141_
rlabel metal3 44072 39032 44072 39032 0 _0142_
rlabel metal2 41160 38836 41160 38836 0 _0143_
rlabel metal2 11032 33208 11032 33208 0 _0144_
rlabel metal2 11256 32592 11256 32592 0 _0145_
rlabel metal3 12264 24584 12264 24584 0 _0146_
rlabel metal2 8904 33600 8904 33600 0 _0147_
rlabel metal2 8120 32424 8120 32424 0 _0148_
rlabel metal2 7896 22008 7896 22008 0 _0149_
rlabel metal2 7560 34272 7560 34272 0 _0150_
rlabel metal3 7000 34216 7000 34216 0 _0151_
rlabel metal2 5600 23800 5600 23800 0 _0152_
rlabel metal2 6328 34104 6328 34104 0 _0153_
rlabel metal2 6328 36008 6328 36008 0 _0154_
rlabel metal2 10136 34440 10136 34440 0 _0155_
rlabel metal2 10248 35672 10248 35672 0 _0156_
rlabel metal2 6776 25592 6776 25592 0 _0157_
rlabel metal2 6888 35952 6888 35952 0 _0158_
rlabel metal2 8120 23576 8120 23576 0 _0159_
rlabel metal2 6888 38024 6888 38024 0 _0160_
rlabel metal2 5880 37352 5880 37352 0 _0161_
rlabel metal2 5320 36176 5320 36176 0 _0162_
rlabel metal2 5712 36680 5712 36680 0 _0163_
rlabel metal2 6888 38528 6888 38528 0 _0164_
rlabel metal2 7280 37352 7280 37352 0 _0165_
rlabel metal2 7056 38808 7056 38808 0 _0166_
rlabel metal2 2800 20104 2800 20104 0 _0167_
rlabel metal2 10024 33544 10024 33544 0 _0168_
rlabel metal2 9688 25480 9688 25480 0 _0169_
rlabel metal2 5768 26880 5768 26880 0 _0170_
rlabel metal3 6776 26264 6776 26264 0 _0171_
rlabel metal2 6328 25536 6328 25536 0 _0172_
rlabel metal3 6272 26488 6272 26488 0 _0173_
rlabel metal2 2968 24696 2968 24696 0 _0174_
rlabel metal2 5320 27552 5320 27552 0 _0175_
rlabel metal3 6440 28056 6440 28056 0 _0176_
rlabel metal3 7000 27272 7000 27272 0 _0177_
rlabel metal2 7112 27832 7112 27832 0 _0178_
rlabel metal2 43848 31528 43848 31528 0 _0179_
rlabel metal2 6440 30968 6440 30968 0 _0180_
rlabel metal2 6776 31192 6776 31192 0 _0181_
rlabel metal2 6440 30464 6440 30464 0 _0182_
rlabel metal3 6608 29400 6608 29400 0 _0183_
rlabel metal2 6216 29680 6216 29680 0 _0184_
rlabel metal2 4984 32200 4984 32200 0 _0185_
rlabel metal2 5992 32144 5992 32144 0 _0186_
rlabel metal2 5768 31472 5768 31472 0 _0187_
rlabel metal3 6776 21448 6776 21448 0 _0188_
rlabel metal2 6720 21000 6720 21000 0 _0189_
rlabel metal2 9016 26936 9016 26936 0 _0190_
rlabel metal2 9016 23912 9016 23912 0 _0191_
rlabel metal3 6608 21672 6608 21672 0 _0192_
rlabel metal2 5768 21952 5768 21952 0 _0193_
rlabel metal2 6216 21056 6216 21056 0 _0194_
rlabel metal2 3080 20328 3080 20328 0 _0195_
rlabel metal2 6104 22064 6104 22064 0 _0196_
rlabel metal2 2968 21896 2968 21896 0 _0197_
rlabel metal2 9520 21784 9520 21784 0 _0198_
rlabel metal3 7896 22232 7896 22232 0 _0199_
rlabel metal3 11760 22232 11760 22232 0 _0200_
rlabel metal2 10696 22848 10696 22848 0 _0201_
rlabel metal2 10584 22792 10584 22792 0 _0202_
rlabel metal3 13384 22456 13384 22456 0 _0203_
rlabel metal2 14056 22624 14056 22624 0 _0204_
rlabel metal2 39704 41832 39704 41832 0 _0205_
rlabel metal3 43820 40488 43820 40488 0 _0206_
rlabel metal2 45360 28056 45360 28056 0 _0207_
rlabel metal2 45192 30688 45192 30688 0 _0208_
rlabel metal2 3640 7056 3640 7056 0 _0209_
rlabel metal3 26264 7392 26264 7392 0 _0210_
rlabel metal2 25928 7728 25928 7728 0 _0211_
rlabel metal2 25368 8456 25368 8456 0 _0212_
rlabel metal3 20384 4872 20384 4872 0 _0213_
rlabel metal2 22232 5488 22232 5488 0 _0214_
rlabel metal2 23016 8288 23016 8288 0 _0215_
rlabel metal3 21000 7448 21000 7448 0 _0216_
rlabel metal2 26712 6272 26712 6272 0 _0217_
rlabel metal2 19544 5544 19544 5544 0 _0218_
rlabel metal2 22456 5152 22456 5152 0 _0219_
rlabel metal2 25032 5376 25032 5376 0 _0220_
rlabel metal2 28168 5376 28168 5376 0 _0221_
rlabel metal2 9576 6664 9576 6664 0 _0222_
rlabel metal2 9296 5992 9296 5992 0 _0223_
rlabel metal3 36736 41160 36736 41160 0 _0224_
rlabel metal2 37688 41048 37688 41048 0 _0225_
rlabel metal2 37128 41552 37128 41552 0 _0226_
rlabel metal2 34216 41216 34216 41216 0 _0227_
rlabel metal2 33880 39984 33880 39984 0 _0228_
rlabel metal2 34104 41440 34104 41440 0 _0229_
rlabel metal2 33768 41552 33768 41552 0 _0230_
rlabel metal3 45360 44296 45360 44296 0 _0231_
rlabel metal2 41272 43456 41272 43456 0 _0232_
rlabel metal2 44856 39200 44856 39200 0 _0233_
rlabel metal2 41720 41272 41720 41272 0 _0234_
rlabel metal2 45248 41160 45248 41160 0 _0235_
rlabel metal2 44576 41160 44576 41160 0 _0236_
rlabel metal2 44072 38752 44072 38752 0 _0237_
rlabel metal3 45640 42056 45640 42056 0 _0238_
rlabel metal2 44968 40096 44968 40096 0 _0239_
rlabel metal2 44744 43876 44744 43876 0 _0240_
rlabel metal2 44800 38808 44800 38808 0 _0241_
rlabel metal2 40152 43876 40152 43876 0 _0242_
rlabel metal2 40656 38808 40656 38808 0 _0243_
rlabel metal2 20552 19488 20552 19488 0 _0244_
rlabel metal2 16856 20440 16856 20440 0 _0245_
rlabel metal2 18312 21392 18312 21392 0 _0246_
rlabel metal3 47432 10584 47432 10584 0 _0247_
rlabel metal3 40712 16072 40712 16072 0 _0248_
rlabel metal2 39480 16128 39480 16128 0 _0249_
rlabel metal2 40152 23184 40152 23184 0 _0250_
rlabel metal2 38920 18144 38920 18144 0 _0251_
rlabel metal2 41272 16632 41272 16632 0 _0252_
rlabel metal2 41552 11368 41552 11368 0 _0253_
rlabel metal2 45192 10808 45192 10808 0 _0254_
rlabel metal3 36960 15848 36960 15848 0 _0255_
rlabel metal2 36456 17248 36456 17248 0 _0256_
rlabel metal2 38472 15120 38472 15120 0 _0257_
rlabel metal2 38864 15960 38864 15960 0 _0258_
rlabel metal3 39536 15960 39536 15960 0 _0259_
rlabel metal2 36120 14224 36120 14224 0 _0260_
rlabel metal3 38724 15400 38724 15400 0 _0261_
rlabel metal2 35672 15624 35672 15624 0 _0262_
rlabel metal2 39256 15008 39256 15008 0 _0263_
rlabel metal2 38024 18312 38024 18312 0 _0264_
rlabel metal2 38080 18536 38080 18536 0 _0265_
rlabel metal2 38696 15708 38696 15708 0 _0266_
rlabel metal2 40824 12992 40824 12992 0 _0267_
rlabel metal2 45080 11312 45080 11312 0 _0268_
rlabel metal2 49448 17584 49448 17584 0 _0269_
rlabel metal2 46312 20328 46312 20328 0 _0270_
rlabel metal2 42168 19544 42168 19544 0 _0271_
rlabel metal3 41216 20776 41216 20776 0 _0272_
rlabel metal2 42168 22008 42168 22008 0 _0273_
rlabel metal2 41832 22680 41832 22680 0 _0274_
rlabel metal2 41944 18760 41944 18760 0 _0275_
rlabel metal3 39816 17640 39816 17640 0 _0276_
rlabel metal2 47432 18088 47432 18088 0 _0277_
rlabel metal2 45640 19376 45640 19376 0 _0278_
rlabel metal2 11928 13832 11928 13832 0 _0279_
rlabel metal2 26488 24920 26488 24920 0 _0280_
rlabel metal2 44856 20048 44856 20048 0 _0281_
rlabel metal2 45528 20216 45528 20216 0 _0282_
rlabel metal2 41496 8568 41496 8568 0 _0283_
rlabel metal2 41888 8120 41888 8120 0 _0284_
rlabel metal2 46536 16296 46536 16296 0 _0285_
rlabel metal2 47096 27160 47096 27160 0 _0286_
rlabel metal3 47208 20104 47208 20104 0 _0287_
rlabel metal2 49112 19432 49112 19432 0 _0288_
rlabel metal3 48328 19768 48328 19768 0 _0289_
rlabel metal2 49784 20048 49784 20048 0 _0290_
rlabel metal2 46984 20160 46984 20160 0 _0291_
rlabel metal2 46592 18536 46592 18536 0 _0292_
rlabel metal2 41608 23184 41608 23184 0 _0293_
rlabel metal2 43512 18256 43512 18256 0 _0294_
rlabel metal2 42952 17248 42952 17248 0 _0295_
rlabel metal3 50232 15960 50232 15960 0 _0296_
rlabel metal2 49224 16688 49224 16688 0 _0297_
rlabel metal2 49560 16464 49560 16464 0 _0298_
rlabel metal2 50120 15596 50120 15596 0 _0299_
rlabel metal3 49504 15960 49504 15960 0 _0300_
rlabel metal2 48776 15624 48776 15624 0 _0301_
rlabel metal2 52920 16128 52920 16128 0 _0302_
rlabel metal3 51800 15960 51800 15960 0 _0303_
rlabel metal2 51800 15624 51800 15624 0 _0304_
rlabel metal3 51744 15176 51744 15176 0 _0305_
rlabel metal2 51576 20384 51576 20384 0 _0306_
rlabel metal2 52024 17584 52024 17584 0 _0307_
rlabel metal2 51240 17920 51240 17920 0 _0308_
rlabel metal3 52192 18424 52192 18424 0 _0309_
rlabel metal2 51352 18200 51352 18200 0 _0310_
rlabel metal3 46536 23800 46536 23800 0 _0311_
rlabel metal2 43848 18032 43848 18032 0 _0312_
rlabel metal2 50120 22624 50120 22624 0 _0313_
rlabel metal2 49784 22232 49784 22232 0 _0314_
rlabel metal2 50008 22008 50008 22008 0 _0315_
rlabel metal3 52080 22232 52080 22232 0 _0316_
rlabel metal3 51128 24808 51128 24808 0 _0317_
rlabel metal2 51688 25760 51688 25760 0 _0318_
rlabel metal2 51912 24920 51912 24920 0 _0319_
rlabel metal2 51520 24920 51520 24920 0 _0320_
rlabel metal2 49112 24976 49112 24976 0 _0321_
rlabel metal2 49224 25760 49224 25760 0 _0322_
rlabel metal2 49560 25312 49560 25312 0 _0323_
rlabel metal2 46984 24696 46984 24696 0 _0324_
rlabel metal2 49784 8960 49784 8960 0 _0325_
rlabel metal2 42392 10640 42392 10640 0 _0326_
rlabel metal2 26040 10304 26040 10304 0 _0327_
rlabel metal2 43960 9296 43960 9296 0 _0328_
rlabel metal2 47880 6552 47880 6552 0 _0329_
rlabel metal2 50008 8400 50008 8400 0 _0330_
rlabel metal2 50680 11200 50680 11200 0 _0331_
rlabel metal2 50456 7112 50456 7112 0 _0332_
rlabel metal2 50120 8568 50120 8568 0 _0333_
rlabel metal2 49784 7000 49784 7000 0 _0334_
rlabel metal3 48384 6552 48384 6552 0 _0335_
rlabel metal2 50568 6496 50568 6496 0 _0336_
rlabel metal2 48888 6608 48888 6608 0 _0337_
rlabel metal2 45192 9408 45192 9408 0 _0338_
rlabel metal2 48552 7112 48552 7112 0 _0339_
rlabel metal3 47096 6664 47096 6664 0 _0340_
rlabel metal2 47656 5432 47656 5432 0 _0341_
rlabel metal2 45976 9016 45976 9016 0 _0342_
rlabel metal3 44240 6664 44240 6664 0 _0343_
rlabel metal3 44688 5208 44688 5208 0 _0344_
rlabel metal2 45136 24024 45136 24024 0 _0345_
rlabel metal2 47152 43400 47152 43400 0 _0346_
rlabel metal2 42000 10472 42000 10472 0 _0347_
rlabel metal2 42840 8680 42840 8680 0 _0348_
rlabel metal3 43960 9016 43960 9016 0 _0349_
rlabel metal2 44968 10584 44968 10584 0 _0350_
rlabel metal2 45752 9464 45752 9464 0 _0351_
rlabel metal2 45192 11872 45192 11872 0 _0352_
rlabel metal2 20272 23240 20272 23240 0 _0353_
rlabel metal2 26544 18312 26544 18312 0 _0354_
rlabel metal2 26264 10696 26264 10696 0 _0355_
rlabel metal2 26712 13104 26712 13104 0 _0356_
rlabel metal2 7448 9856 7448 9856 0 _0357_
rlabel metal2 27608 18704 27608 18704 0 _0358_
rlabel metal2 31864 10920 31864 10920 0 _0359_
rlabel metal3 40208 10024 40208 10024 0 _0360_
rlabel metal2 38808 10640 38808 10640 0 _0361_
rlabel metal2 33432 10136 33432 10136 0 _0362_
rlabel metal3 32424 8792 32424 8792 0 _0363_
rlabel metal2 34328 12544 34328 12544 0 _0364_
rlabel metal3 38668 12376 38668 12376 0 _0365_
rlabel metal2 39032 12152 39032 12152 0 _0366_
rlabel metal2 32200 11648 32200 11648 0 _0367_
rlabel metal2 32536 11760 32536 11760 0 _0368_
rlabel metal2 43848 23800 43848 23800 0 _0369_
rlabel metal2 31752 11704 31752 11704 0 _0370_
rlabel metal2 35896 12600 35896 12600 0 _0371_
rlabel metal2 36120 12600 36120 12600 0 _0372_
rlabel metal2 26712 21952 26712 21952 0 _0373_
rlabel metal2 39256 7952 39256 7952 0 _0374_
rlabel metal3 38192 13720 38192 13720 0 _0375_
rlabel metal2 40040 14168 40040 14168 0 _0376_
rlabel metal2 50176 23912 50176 23912 0 _0377_
rlabel metal2 38808 12544 38808 12544 0 _0378_
rlabel metal3 40040 12824 40040 12824 0 _0379_
rlabel metal2 41048 12992 41048 12992 0 _0380_
rlabel metal2 36624 9016 36624 9016 0 _0381_
rlabel metal2 36232 9968 36232 9968 0 _0382_
rlabel metal3 37016 9128 37016 9128 0 _0383_
rlabel metal2 34776 8456 34776 8456 0 _0384_
rlabel metal3 35392 8120 35392 8120 0 _0385_
rlabel metal2 36680 8120 36680 8120 0 _0386_
rlabel metal2 38920 8316 38920 8316 0 _0387_
rlabel metal2 38360 8064 38360 8064 0 _0388_
rlabel metal3 37520 7448 37520 7448 0 _0389_
rlabel metal2 19936 18984 19936 18984 0 _0390_
rlabel metal2 23800 8344 23800 8344 0 _0391_
rlabel metal2 39088 6888 39088 6888 0 _0392_
rlabel metal2 39368 7896 39368 7896 0 _0393_
rlabel metal2 40712 8456 40712 8456 0 _0394_
rlabel metal2 24136 6272 24136 6272 0 _0395_
rlabel metal2 26040 8176 26040 8176 0 _0396_
rlabel metal2 40936 7112 40936 7112 0 _0397_
rlabel metal2 40824 7336 40824 7336 0 _0398_
rlabel metal2 26320 9240 26320 9240 0 _0399_
rlabel metal3 28168 11368 28168 11368 0 _0400_
rlabel metal2 26376 13104 26376 13104 0 _0401_
rlabel metal2 24472 16016 24472 16016 0 _0402_
rlabel metal2 24360 17248 24360 17248 0 _0403_
rlabel metal2 26376 14000 26376 14000 0 _0404_
rlabel metal3 24080 12152 24080 12152 0 _0405_
rlabel metal2 24080 12264 24080 12264 0 _0406_
rlabel metal3 24752 10696 24752 10696 0 _0407_
rlabel metal2 25312 15960 25312 15960 0 _0408_
rlabel metal2 25592 16072 25592 16072 0 _0409_
rlabel metal2 23128 17528 23128 17528 0 _0410_
rlabel metal2 23240 13776 23240 13776 0 _0411_
rlabel metal2 23688 16184 23688 16184 0 _0412_
rlabel metal2 23520 19656 23520 19656 0 _0413_
rlabel metal2 23912 21056 23912 21056 0 _0414_
rlabel metal2 23912 11284 23912 11284 0 _0415_
rlabel metal2 23800 19600 23800 19600 0 _0416_
rlabel metal2 27608 22008 27608 22008 0 _0417_
rlabel metal2 27216 21784 27216 21784 0 _0418_
rlabel metal2 11704 39200 11704 39200 0 _0419_
rlabel metal2 26264 46200 26264 46200 0 _0420_
rlabel metal2 45976 47600 45976 47600 0 _0421_
rlabel metal2 33544 8568 33544 8568 0 _0422_
rlabel metal2 32312 5432 32312 5432 0 _0423_
rlabel metal2 43736 25200 43736 25200 0 _0424_
rlabel metal2 29176 26096 29176 26096 0 _0425_
rlabel metal2 43960 22344 43960 22344 0 _0426_
rlabel metal2 39312 23016 39312 23016 0 _0427_
rlabel metal2 31864 27160 31864 27160 0 _0428_
rlabel metal2 30520 31304 30520 31304 0 _0429_
rlabel metal2 31472 26824 31472 26824 0 _0430_
rlabel metal2 36232 44856 36232 44856 0 _0431_
rlabel metal2 34440 24360 34440 24360 0 _0432_
rlabel metal2 30856 27272 30856 27272 0 _0433_
rlabel metal2 33880 17472 33880 17472 0 _0434_
rlabel metal2 14616 13216 14616 13216 0 _0435_
rlabel metal3 39844 21336 39844 21336 0 _0436_
rlabel metal2 34216 30296 34216 30296 0 _0437_
rlabel metal2 31080 31360 31080 31360 0 _0438_
rlabel metal2 31584 31976 31584 31976 0 _0439_
rlabel metal2 44632 17808 44632 17808 0 _0440_
rlabel metal2 31528 30016 31528 30016 0 _0441_
rlabel metal2 31192 29624 31192 29624 0 _0442_
rlabel metal2 34888 32872 34888 32872 0 _0443_
rlabel metal3 41496 18424 41496 18424 0 _0444_
rlabel metal2 34496 31192 34496 31192 0 _0445_
rlabel metal2 33992 34328 33992 34328 0 _0446_
rlabel metal2 33936 31752 33936 31752 0 _0447_
rlabel metal3 20104 16744 20104 16744 0 _0448_
rlabel metal2 34048 31192 34048 31192 0 _0449_
rlabel metal2 33656 34608 33656 34608 0 _0450_
rlabel metal3 16744 17416 16744 17416 0 _0451_
rlabel metal2 34720 27608 34720 27608 0 _0452_
rlabel metal2 34328 34552 34328 34552 0 _0453_
rlabel metal2 15904 17080 15904 17080 0 _0454_
rlabel metal2 35224 30016 35224 30016 0 _0455_
rlabel metal2 34832 34776 34832 34776 0 _0456_
rlabel metal2 49056 15624 49056 15624 0 _0457_
rlabel metal3 49112 33320 49112 33320 0 _0458_
rlabel metal2 49448 34888 49448 34888 0 _0459_
rlabel metal2 38808 35728 38808 35728 0 _0460_
rlabel metal2 42168 23464 42168 23464 0 _0461_
rlabel metal2 42504 25900 42504 25900 0 _0462_
rlabel metal3 39872 36456 39872 36456 0 _0463_
rlabel metal2 43736 33936 43736 33936 0 _0464_
rlabel metal2 43568 23352 43568 23352 0 _0465_
rlabel metal2 40824 24640 40824 24640 0 _0466_
rlabel metal2 42168 30632 42168 30632 0 _0467_
rlabel metal2 43624 31416 43624 31416 0 _0468_
rlabel metal2 43960 32480 43960 32480 0 _0469_
rlabel metal2 45080 32928 45080 32928 0 _0470_
rlabel metal2 42056 20552 42056 20552 0 _0471_
rlabel metal2 30408 21784 30408 21784 0 _0472_
rlabel metal2 30016 22456 30016 22456 0 _0473_
rlabel metal2 33544 20664 33544 20664 0 _0474_
rlabel metal2 40600 21448 40600 21448 0 _0475_
rlabel metal3 40824 24696 40824 24696 0 _0476_
rlabel metal2 39816 24024 39816 24024 0 _0477_
rlabel metal3 44184 21504 44184 21504 0 _0478_
rlabel metal3 46984 32312 46984 32312 0 _0479_
rlabel metal2 50176 31976 50176 31976 0 _0480_
rlabel metal2 41608 34832 41608 34832 0 _0481_
rlabel metal3 42784 34888 42784 34888 0 _0482_
rlabel metal2 38024 21560 38024 21560 0 _0483_
rlabel metal2 41216 35672 41216 35672 0 _0484_
rlabel metal2 31192 21616 31192 21616 0 _0485_
rlabel metal2 39144 22624 39144 22624 0 _0486_
rlabel metal3 44408 22120 44408 22120 0 _0487_
rlabel metal2 49448 48440 49448 48440 0 _0488_
rlabel metal3 47656 34776 47656 34776 0 _0489_
rlabel metal2 31752 35672 31752 35672 0 _0490_
rlabel metal2 37128 19936 37128 19936 0 _0491_
rlabel metal2 37520 20104 37520 20104 0 _0492_
rlabel metal2 44128 25368 44128 25368 0 _0493_
rlabel metal2 46200 36792 46200 36792 0 _0494_
rlabel metal3 50568 44072 50568 44072 0 _0495_
rlabel metal2 42280 33544 42280 33544 0 _0496_
rlabel metal2 24136 30576 24136 30576 0 _0497_
rlabel metal2 42056 32312 42056 32312 0 _0498_
rlabel metal3 40236 32536 40236 32536 0 _0499_
rlabel metal2 42616 33208 42616 33208 0 _0500_
rlabel metal2 50904 33768 50904 33768 0 _0501_
rlabel metal2 42728 33992 42728 33992 0 _0502_
rlabel metal2 23800 29736 23800 29736 0 _0503_
rlabel metal2 24808 31808 24808 31808 0 _0504_
rlabel metal2 39032 34888 39032 34888 0 _0505_
rlabel metal2 39256 32816 39256 32816 0 _0506_
rlabel metal2 47208 34888 47208 34888 0 _0507_
rlabel metal2 50904 35448 50904 35448 0 _0508_
rlabel metal2 48552 42168 48552 42168 0 _0509_
rlabel metal2 51912 43960 51912 43960 0 _0510_
rlabel metal2 43848 34608 43848 34608 0 _0511_
rlabel metal2 24360 32032 24360 32032 0 _0512_
rlabel metal3 41384 34104 41384 34104 0 _0513_
rlabel metal2 49056 39144 49056 39144 0 _0514_
rlabel metal2 49896 42280 49896 42280 0 _0515_
rlabel metal2 44184 36064 44184 36064 0 _0516_
rlabel metal2 25032 31752 25032 31752 0 _0517_
rlabel metal2 40152 35168 40152 35168 0 _0518_
rlabel metal3 46872 37688 46872 37688 0 _0519_
rlabel metal2 49896 39256 49896 39256 0 _0520_
rlabel metal2 41720 35952 41720 35952 0 _0521_
rlabel metal2 40376 33376 40376 33376 0 _0522_
rlabel metal2 39256 34664 39256 34664 0 _0523_
rlabel metal3 47320 43736 47320 43736 0 _0524_
rlabel metal2 51464 44296 51464 44296 0 _0525_
rlabel metal2 33712 44296 33712 44296 0 _0526_
rlabel metal2 19320 34440 19320 34440 0 _0527_
rlabel metal2 19880 35224 19880 35224 0 _0528_
rlabel metal2 18592 35560 18592 35560 0 _0529_
rlabel metal2 18536 35056 18536 35056 0 _0530_
rlabel metal2 18984 36680 18984 36680 0 _0531_
rlabel metal2 18200 36568 18200 36568 0 _0532_
rlabel metal2 18312 36792 18312 36792 0 _0533_
rlabel metal2 16856 36792 16856 36792 0 _0534_
rlabel metal2 16576 36344 16576 36344 0 _0535_
rlabel metal2 17976 36904 17976 36904 0 _0536_
rlabel metal2 18928 41384 18928 41384 0 _0537_
rlabel metal2 29288 37688 29288 37688 0 _0538_
rlabel metal3 29064 38024 29064 38024 0 _0539_
rlabel metal3 29176 38248 29176 38248 0 _0540_
rlabel metal3 28896 38360 28896 38360 0 _0541_
rlabel metal2 29176 38584 29176 38584 0 _0542_
rlabel metal2 26264 36064 26264 36064 0 _0543_
rlabel metal2 22904 36120 22904 36120 0 _0544_
rlabel metal2 24304 36568 24304 36568 0 _0545_
rlabel metal3 23520 36344 23520 36344 0 _0546_
rlabel metal2 25704 37016 25704 37016 0 _0547_
rlabel metal2 31976 42560 31976 42560 0 _0548_
rlabel metal2 47544 44912 47544 44912 0 _0549_
rlabel metal2 47768 47712 47768 47712 0 _0550_
rlabel metal2 34160 44296 34160 44296 0 _0551_
rlabel metal2 38864 44520 38864 44520 0 _0552_
rlabel metal2 47768 46480 47768 46480 0 _0553_
rlabel metal2 46816 48328 46816 48328 0 _0554_
rlabel metal3 49392 47544 49392 47544 0 _0555_
rlabel metal2 50624 47320 50624 47320 0 _0556_
rlabel metal2 49784 50288 49784 50288 0 _0557_
rlabel metal2 50008 50232 50008 50232 0 _0558_
rlabel metal2 49896 50680 49896 50680 0 _0559_
rlabel metal3 48328 45304 48328 45304 0 _0560_
rlabel metal2 48216 46256 48216 46256 0 _0561_
rlabel metal2 48272 45192 48272 45192 0 _0562_
rlabel metal2 48104 45640 48104 45640 0 _0563_
rlabel metal2 47544 45752 47544 45752 0 _0564_
rlabel metal2 47600 43736 47600 43736 0 _0565_
rlabel metal2 45752 27552 45752 27552 0 _0566_
rlabel metal2 46760 28280 46760 28280 0 _0567_
rlabel metal2 47432 28952 47432 28952 0 _0568_
rlabel metal2 47656 29512 47656 29512 0 _0569_
rlabel metal2 25928 25872 25928 25872 0 _0570_
rlabel metal2 26152 25088 26152 25088 0 _0571_
rlabel metal2 26768 24472 26768 24472 0 _0572_
rlabel metal2 29512 24696 29512 24696 0 _0573_
rlabel metal2 27384 31416 27384 31416 0 _0574_
rlabel metal2 25704 28616 25704 28616 0 _0575_
rlabel metal2 22680 31808 22680 31808 0 _0576_
rlabel metal2 26824 31752 26824 31752 0 _0577_
rlabel metal2 26208 30184 26208 30184 0 _0578_
rlabel metal2 25816 32592 25816 32592 0 _0579_
rlabel metal2 24192 26488 24192 26488 0 _0580_
rlabel metal3 22064 30184 22064 30184 0 _0581_
rlabel metal3 21952 30968 21952 30968 0 _0582_
rlabel metal2 22456 33768 22456 33768 0 _0583_
rlabel metal2 22008 30968 22008 30968 0 _0584_
rlabel metal2 21672 33040 21672 33040 0 _0585_
rlabel metal2 21672 26992 21672 26992 0 _0586_
rlabel metal2 21504 27048 21504 27048 0 _0587_
rlabel metal2 23688 28056 23688 28056 0 _0588_
rlabel metal2 23128 28168 23128 28168 0 _0589_
rlabel metal2 39144 26992 39144 26992 0 _0590_
rlabel metal2 39704 25704 39704 25704 0 _0591_
rlabel metal2 39368 28112 39368 28112 0 _0592_
rlabel metal2 34608 23912 34608 23912 0 _0593_
rlabel metal3 36456 23800 36456 23800 0 _0594_
rlabel metal2 40040 27832 40040 27832 0 _0595_
rlabel metal3 34104 19208 34104 19208 0 _0596_
rlabel metal2 33992 18312 33992 18312 0 _0597_
rlabel metal3 31864 18424 31864 18424 0 _0598_
rlabel metal2 40488 29008 40488 29008 0 _0599_
rlabel metal2 40824 29120 40824 29120 0 _0600_
rlabel metal2 26264 39704 26264 39704 0 _0601_
rlabel metal3 36904 28616 36904 28616 0 _0602_
rlabel metal2 37688 28616 37688 28616 0 _0603_
rlabel metal2 40208 26824 40208 26824 0 _0604_
rlabel metal2 40432 28056 40432 28056 0 _0605_
rlabel metal2 39704 29008 39704 29008 0 _0606_
rlabel metal3 32200 47208 32200 47208 0 _0607_
rlabel metal3 24864 42616 24864 42616 0 _0608_
rlabel metal2 14504 44240 14504 44240 0 _0609_
rlabel metal2 11256 42112 11256 42112 0 _0610_
rlabel metal3 36792 44184 36792 44184 0 _0611_
rlabel metal2 38808 43736 38808 43736 0 _0612_
rlabel metal2 14840 45528 14840 45528 0 _0613_
rlabel metal3 24024 45640 24024 45640 0 _0614_
rlabel metal3 24360 42728 24360 42728 0 _0615_
rlabel metal3 25928 42840 25928 42840 0 _0616_
rlabel metal2 21560 40824 21560 40824 0 _0617_
rlabel metal2 25648 39592 25648 39592 0 _0618_
rlabel metal2 24696 42336 24696 42336 0 _0619_
rlabel metal2 34552 44800 34552 44800 0 _0620_
rlabel metal2 22792 43344 22792 43344 0 _0621_
rlabel metal3 22456 49056 22456 49056 0 _0622_
rlabel metal2 25256 40264 25256 40264 0 _0623_
rlabel metal2 24024 39592 24024 39592 0 _0624_
rlabel metal2 14728 44016 14728 44016 0 _0625_
rlabel metal3 20720 41048 20720 41048 0 _0626_
rlabel metal3 13216 41160 13216 41160 0 _0627_
rlabel metal2 20552 41216 20552 41216 0 _0628_
rlabel metal2 22904 41328 22904 41328 0 _0629_
rlabel metal2 19208 40824 19208 40824 0 _0630_
rlabel metal3 18312 41048 18312 41048 0 _0631_
rlabel metal2 12152 42056 12152 42056 0 _0632_
rlabel metal2 21784 43512 21784 43512 0 _0633_
rlabel metal2 21336 43176 21336 43176 0 _0634_
rlabel metal2 18312 41832 18312 41832 0 _0635_
rlabel metal2 6888 12768 6888 12768 0 _0636_
rlabel metal2 22176 45080 22176 45080 0 _0637_
rlabel metal3 23520 50456 23520 50456 0 _0638_
rlabel metal3 24976 48888 24976 48888 0 _0639_
rlabel metal2 23016 49392 23016 49392 0 _0640_
rlabel metal2 21392 49560 21392 49560 0 _0641_
rlabel metal2 19880 49840 19880 49840 0 _0642_
rlabel metal2 20888 50568 20888 50568 0 _0643_
rlabel metal3 23912 47320 23912 47320 0 _0644_
rlabel metal3 23688 48776 23688 48776 0 _0645_
rlabel metal2 22344 49112 22344 49112 0 _0646_
rlabel metal2 22792 48216 22792 48216 0 _0647_
rlabel metal2 23576 50120 23576 50120 0 _0648_
rlabel metal2 25704 49504 25704 49504 0 _0649_
rlabel metal2 26488 50484 26488 50484 0 _0650_
rlabel metal2 23240 50064 23240 50064 0 _0651_
rlabel metal2 26152 50624 26152 50624 0 _0652_
rlabel metal3 27272 49784 27272 49784 0 _0653_
rlabel metal2 25928 48496 25928 48496 0 _0654_
rlabel metal2 26488 49448 26488 49448 0 _0655_
rlabel via2 25144 44968 25144 44968 0 _0656_
rlabel metal2 22344 44800 22344 44800 0 _0657_
rlabel metal2 22680 45528 22680 45528 0 _0658_
rlabel metal3 21000 46088 21000 46088 0 _0659_
rlabel metal2 23128 45472 23128 45472 0 _0660_
rlabel metal3 21952 46648 21952 46648 0 _0661_
rlabel metal3 24416 44520 24416 44520 0 _0662_
rlabel metal2 19992 44744 19992 44744 0 _0663_
rlabel metal2 20552 46368 20552 46368 0 _0664_
rlabel metal2 21000 47040 21000 47040 0 _0665_
rlabel metal2 21056 47432 21056 47432 0 _0666_
rlabel metal3 18312 44296 18312 44296 0 _0667_
rlabel metal2 16520 43792 16520 43792 0 _0668_
rlabel metal2 16744 44968 16744 44968 0 _0669_
rlabel metal2 16184 45360 16184 45360 0 _0670_
rlabel metal2 17416 46144 17416 46144 0 _0671_
rlabel metal2 16632 45864 16632 45864 0 _0672_
rlabel metal2 16296 46144 16296 46144 0 _0673_
rlabel metal3 21952 44856 21952 44856 0 _0674_
rlabel metal2 13384 44744 13384 44744 0 _0675_
rlabel metal3 12600 45192 12600 45192 0 _0676_
rlabel metal2 11816 44408 11816 44408 0 _0677_
rlabel metal3 10752 43848 10752 43848 0 _0678_
rlabel metal3 10248 44072 10248 44072 0 _0679_
rlabel metal2 11256 40040 11256 40040 0 _0680_
rlabel metal2 10416 45752 10416 45752 0 _0681_
rlabel metal2 11032 45360 11032 45360 0 _0682_
rlabel metal3 13384 45080 13384 45080 0 _0683_
rlabel metal2 12376 45080 12376 45080 0 _0684_
rlabel metal2 12152 41440 12152 41440 0 _0685_
rlabel metal2 12152 43876 12152 43876 0 _0686_
rlabel metal2 12712 42224 12712 42224 0 _0687_
rlabel metal2 13440 41944 13440 41944 0 _0688_
rlabel metal3 11704 41944 11704 41944 0 _0689_
rlabel metal2 10920 42000 10920 42000 0 _0690_
rlabel metal2 14560 39816 14560 39816 0 _0691_
rlabel metal2 13384 39480 13384 39480 0 _0692_
rlabel metal2 13944 40376 13944 40376 0 _0693_
rlabel metal2 13944 9856 13944 9856 0 _0694_
rlabel metal2 49112 45640 49112 45640 0 _0695_
rlabel metal3 37072 46200 37072 46200 0 _0696_
rlabel metal2 39256 47936 39256 47936 0 _0697_
rlabel metal2 39032 49112 39032 49112 0 _0698_
rlabel metal2 39256 45584 39256 45584 0 _0699_
rlabel metal2 34888 49112 34888 49112 0 _0700_
rlabel metal2 33432 47432 33432 47432 0 _0701_
rlabel metal2 42056 49840 42056 49840 0 _0702_
rlabel metal2 34328 49560 34328 49560 0 _0703_
rlabel metal3 37240 49672 37240 49672 0 _0704_
rlabel metal2 39480 47376 39480 47376 0 _0705_
rlabel metal3 40432 49672 40432 49672 0 _0706_
rlabel metal2 42504 47936 42504 47936 0 _0707_
rlabel metal2 42952 46704 42952 46704 0 _0708_
rlabel metal2 42728 46200 42728 46200 0 _0709_
rlabel metal2 42280 45808 42280 45808 0 _0710_
rlabel metal2 37016 46200 37016 46200 0 _0711_
rlabel metal2 39928 43008 39928 43008 0 _0712_
rlabel metal3 40096 44072 40096 44072 0 _0713_
rlabel metal2 34552 42392 34552 42392 0 _0714_
rlabel metal3 15680 22568 15680 22568 0 _0715_
rlabel metal2 16184 30912 16184 30912 0 _0716_
rlabel metal2 16520 30912 16520 30912 0 _0717_
rlabel metal3 15232 32648 15232 32648 0 _0718_
rlabel metal2 15176 34104 15176 34104 0 _0719_
rlabel metal2 15064 32088 15064 32088 0 _0720_
rlabel metal2 15512 33656 15512 33656 0 _0721_
rlabel metal3 13888 34104 13888 34104 0 _0722_
rlabel metal2 13552 35560 13552 35560 0 _0723_
rlabel metal2 12264 34888 12264 34888 0 _0724_
rlabel metal2 15624 32816 15624 32816 0 _0725_
rlabel metal3 12544 17752 12544 17752 0 _0726_
rlabel metal2 8344 14616 8344 14616 0 _0727_
rlabel metal2 19768 28000 19768 28000 0 _0728_
rlabel metal2 20384 28728 20384 28728 0 _0729_
rlabel metal2 18312 28840 18312 28840 0 _0730_
rlabel metal2 18424 29568 18424 29568 0 _0731_
rlabel metal2 18536 25900 18536 25900 0 _0732_
rlabel metal2 19152 24024 19152 24024 0 _0733_
rlabel metal2 19096 30072 19096 30072 0 _0734_
rlabel metal3 19096 25480 19096 25480 0 _0735_
rlabel metal3 19040 25704 19040 25704 0 _0736_
rlabel metal2 18704 24808 18704 24808 0 _0737_
rlabel metal2 16744 22680 16744 22680 0 _0738_
rlabel metal2 6440 14896 6440 14896 0 _0739_
rlabel metal2 5768 11928 5768 11928 0 _0740_
rlabel metal2 32088 19992 32088 19992 0 _0741_
rlabel metal3 9464 14616 9464 14616 0 _0742_
rlabel metal2 8792 14504 8792 14504 0 _0743_
rlabel metal2 8904 14056 8904 14056 0 _0744_
rlabel metal2 6104 13944 6104 13944 0 _0745_
rlabel metal2 6216 14448 6216 14448 0 _0746_
rlabel metal3 8568 17640 8568 17640 0 _0747_
rlabel metal2 8232 19880 8232 19880 0 _0748_
rlabel metal2 10136 19992 10136 19992 0 _0749_
rlabel metal2 8680 18648 8680 18648 0 _0750_
rlabel metal2 8176 12712 8176 12712 0 _0751_
rlabel metal3 5432 12936 5432 12936 0 _0752_
rlabel metal2 6440 12040 6440 12040 0 _0753_
rlabel metal3 23464 20104 23464 20104 0 _0754_
rlabel metal2 12712 14224 12712 14224 0 _0755_
rlabel metal2 9184 11592 9184 11592 0 _0756_
rlabel metal2 6776 14280 6776 14280 0 _0757_
rlabel metal2 6664 13048 6664 13048 0 _0758_
rlabel metal2 7448 12376 7448 12376 0 _0759_
rlabel metal3 7448 12096 7448 12096 0 _0760_
rlabel metal2 5992 15680 5992 15680 0 _0761_
rlabel metal2 6384 15512 6384 15512 0 _0762_
rlabel metal2 6328 10920 6328 10920 0 _0763_
rlabel metal2 6104 16520 6104 16520 0 _0764_
rlabel metal2 5936 10584 5936 10584 0 _0765_
rlabel metal2 6664 10864 6664 10864 0 _0766_
rlabel metal2 13608 15624 13608 15624 0 _0767_
rlabel metal2 11480 13384 11480 13384 0 _0768_
rlabel metal3 10920 10584 10920 10584 0 _0769_
rlabel metal2 10192 10808 10192 10808 0 _0770_
rlabel metal2 8792 7224 8792 7224 0 _0771_
rlabel metal3 10248 11592 10248 11592 0 _0772_
rlabel metal2 9576 10920 9576 10920 0 _0773_
rlabel metal2 11592 9856 11592 9856 0 _0774_
rlabel metal3 13720 9800 13720 9800 0 _0775_
rlabel metal2 11480 11872 11480 11872 0 _0776_
rlabel metal2 11256 10584 11256 10584 0 _0777_
rlabel metal3 13720 9688 13720 9688 0 _0778_
rlabel metal2 14952 13216 14952 13216 0 _0779_
rlabel metal3 13160 11368 13160 11368 0 _0780_
rlabel metal2 12488 10248 12488 10248 0 _0781_
rlabel metal2 14280 9632 14280 9632 0 _0782_
rlabel metal2 17640 13832 17640 13832 0 _0783_
rlabel metal2 13608 11312 13608 11312 0 _0784_
rlabel metal2 14112 10024 14112 10024 0 _0785_
rlabel metal2 18648 11872 18648 11872 0 _0786_
rlabel metal2 16016 16856 16016 16856 0 _0787_
rlabel metal2 15400 12040 15400 12040 0 _0788_
rlabel metal2 16016 12152 16016 12152 0 _0789_
rlabel metal2 17976 16968 17976 16968 0 _0790_
rlabel metal2 18536 13888 18536 13888 0 _0791_
rlabel metal2 17416 16912 17416 16912 0 _0792_
rlabel metal2 15736 16016 15736 16016 0 _0793_
rlabel metal3 18144 12936 18144 12936 0 _0794_
rlabel metal2 17808 12152 17808 12152 0 _0795_
rlabel metal2 17528 16408 17528 16408 0 _0796_
rlabel metal2 17752 14448 17752 14448 0 _0797_
rlabel metal2 17920 14280 17920 14280 0 _0798_
rlabel metal2 15512 16856 15512 16856 0 _0799_
rlabel metal2 17416 16240 17416 16240 0 _0800_
rlabel metal3 17024 16744 17024 16744 0 _0801_
rlabel metal2 12936 15624 12936 15624 0 _0802_
rlabel metal2 15400 16576 15400 16576 0 _0803_
rlabel metal3 14056 16856 14056 16856 0 _0804_
rlabel metal3 12152 16856 12152 16856 0 _0805_
rlabel metal2 10360 27496 10360 27496 0 _0806_
rlabel metal2 7560 18760 7560 18760 0 _0807_
rlabel metal2 11816 22848 11816 22848 0 _0808_
rlabel metal2 11928 26152 11928 26152 0 _0809_
rlabel metal2 5600 21560 5600 21560 0 _0810_
rlabel metal2 6832 26264 6832 26264 0 _0811_
rlabel metal2 9912 29344 9912 29344 0 _0812_
rlabel metal3 11816 29288 11816 29288 0 _0813_
rlabel metal3 9968 28728 9968 28728 0 _0814_
rlabel metal2 10024 30296 10024 30296 0 _0815_
rlabel metal2 9968 28840 9968 28840 0 _0816_
rlabel metal2 9576 22624 9576 22624 0 _0817_
rlabel metal2 9800 34888 9800 34888 0 _0818_
rlabel metal2 9912 30688 9912 30688 0 _0819_
rlabel metal3 7476 38808 7476 38808 0 _0820_
rlabel metal3 12040 26544 12040 26544 0 _0821_
rlabel metal2 11592 26096 11592 26096 0 _0822_
rlabel metal3 11032 25368 11032 25368 0 _0823_
rlabel metal2 12600 26376 12600 26376 0 _0824_
rlabel metal2 11256 26544 11256 26544 0 _0825_
rlabel metal3 13104 24696 13104 24696 0 _0826_
rlabel metal2 53256 3304 53256 3304 0 addr[0]
rlabel metal2 53312 6440 53312 6440 0 addr[1]
rlabel metal2 53368 7952 53368 7952 0 addr[2]
rlabel metal2 42952 2184 42952 2184 0 bus_cyc
rlabel metal2 47544 2058 47544 2058 0 bus_we
rlabel metal2 46648 45192 46648 45192 0 clknet_0_wb_clk_i
rlabel metal3 6440 8232 6440 8232 0 clknet_4_0_0_wb_clk_i
rlabel metal2 51464 13832 51464 13832 0 clknet_4_10_0_wb_clk_i
rlabel metal2 47992 22736 47992 22736 0 clknet_4_11_0_wb_clk_i
rlabel metal2 39256 39480 39256 39480 0 clknet_4_12_0_wb_clk_i
rlabel metal2 32256 50568 32256 50568 0 clknet_4_13_0_wb_clk_i
rlabel metal2 50176 44968 50176 44968 0 clknet_4_14_0_wb_clk_i
rlabel metal2 50456 46872 50456 46872 0 clknet_4_15_0_wb_clk_i
rlabel metal2 4872 11928 4872 11928 0 clknet_4_1_0_wb_clk_i
rlabel metal3 25648 13720 25648 13720 0 clknet_4_2_0_wb_clk_i
rlabel metal3 20496 15288 20496 15288 0 clknet_4_3_0_wb_clk_i
rlabel metal2 1736 21280 1736 21280 0 clknet_4_4_0_wb_clk_i
rlabel metal2 7112 44296 7112 44296 0 clknet_4_5_0_wb_clk_i
rlabel metal2 16912 21784 16912 21784 0 clknet_4_6_0_wb_clk_i
rlabel metal2 13048 47040 13048 47040 0 clknet_4_7_0_wb_clk_i
rlabel metal2 44184 16016 44184 16016 0 clknet_4_8_0_wb_clk_i
rlabel metal2 38808 24360 38808 24360 0 clknet_4_9_0_wb_clk_i
rlabel metal3 53746 11256 53746 11256 0 data_in[0]
rlabel metal3 53802 13944 53802 13944 0 data_in[1]
rlabel metal3 53256 16744 53256 16744 0 data_in[2]
rlabel metal2 53256 19264 53256 19264 0 data_in[3]
rlabel metal2 53256 21840 53256 21840 0 data_in[4]
rlabel metal3 53746 24696 53746 24696 0 data_in[5]
rlabel metal3 53802 27384 53802 27384 0 data_in[6]
rlabel metal3 53746 30072 53746 30072 0 data_in[7]
rlabel metal2 53032 33320 53032 33320 0 data_out[0]
rlabel metal2 53032 36232 53032 36232 0 data_out[1]
rlabel metal3 53634 38136 53634 38136 0 data_out[2]
rlabel metal2 51912 41048 51912 41048 0 data_out[3]
rlabel metal2 53032 43456 53032 43456 0 data_out[4]
rlabel metal2 53032 47096 53032 47096 0 data_out[5]
rlabel metal2 51912 49000 51912 49000 0 data_out[6]
rlabel metal3 52682 51576 52682 51576 0 data_out[7]
rlabel metal2 2744 2086 2744 2086 0 io_in
rlabel metal2 7224 2086 7224 2086 0 io_out[0]
rlabel metal2 11704 2422 11704 2422 0 io_out[1]
rlabel metal2 52024 2198 52024 2198 0 irq3
rlabel metal2 39480 44688 39480 44688 0 net1
rlabel metal2 45192 18088 45192 18088 0 net10
rlabel metal2 51240 17584 51240 17584 0 net11
rlabel metal2 49784 23520 49784 23520 0 net12
rlabel metal3 47544 26376 47544 26376 0 net13
rlabel metal2 49224 26684 49224 26684 0 net14
rlabel metal2 3304 5376 3304 5376 0 net15
rlabel metal2 41832 51240 41832 51240 0 net16
rlabel metal2 10584 5824 10584 5824 0 net17
rlabel metal2 49560 33264 49560 33264 0 net18
rlabel metal2 49784 35616 49784 35616 0 net19
rlabel metal2 52696 4312 52696 4312 0 net2
rlabel metal2 49672 38416 49672 38416 0 net20
rlabel metal2 50120 41160 50120 41160 0 net21
rlabel metal2 51184 43512 51184 43512 0 net22
rlabel metal2 50680 45976 50680 45976 0 net23
rlabel metal2 49728 45752 49728 45752 0 net24
rlabel metal3 52640 44968 52640 44968 0 net25
rlabel metal2 11928 3472 11928 3472 0 net26
rlabel metal2 14392 4424 14392 4424 0 net27
rlabel metal2 53256 4032 53256 4032 0 net28
rlabel metal2 20664 2030 20664 2030 0 net29
rlabel metal3 52136 6664 52136 6664 0 net3
rlabel metal2 25256 4424 25256 4424 0 net30
rlabel metal2 16184 2030 16184 2030 0 net31
rlabel metal2 29624 2058 29624 2058 0 net32
rlabel metal2 52920 8260 52920 8260 0 net4
rlabel metal2 44352 24584 44352 24584 0 net5
rlabel metal2 44856 24528 44856 24528 0 net6
rlabel metal2 52920 12768 52920 12768 0 net7
rlabel metal2 52696 14840 52696 14840 0 net8
rlabel metal3 47208 16968 47208 16968 0 net9
rlabel metal2 41272 52906 41272 52906 0 rst
rlabel metal2 41608 19656 41608 19656 0 spi.busy
rlabel metal2 52808 9744 52808 9744 0 spi.counter\[0\]
rlabel metal2 52752 7448 52752 7448 0 spi.counter\[1\]
rlabel metal2 49224 6440 49224 6440 0 spi.counter\[2\]
rlabel metal2 46536 5152 46536 5152 0 spi.counter\[3\]
rlabel metal3 48608 9688 48608 9688 0 spi.counter\[4\]
rlabel metal2 26152 8848 26152 8848 0 spi.data_in_buff\[0\]
rlabel metal3 24752 12712 24752 12712 0 spi.data_in_buff\[1\]
rlabel metal3 24080 8120 24080 8120 0 spi.data_in_buff\[2\]
rlabel metal2 23520 7560 23520 7560 0 spi.data_in_buff\[3\]
rlabel metal2 22792 7280 22792 7280 0 spi.data_in_buff\[4\]
rlabel metal3 23968 6104 23968 6104 0 spi.data_in_buff\[5\]
rlabel metal2 24584 6664 24584 6664 0 spi.data_in_buff\[6\]
rlabel metal2 27384 7728 27384 7728 0 spi.data_in_buff\[7\]
rlabel metal2 46760 20888 46760 20888 0 spi.data_out_buff\[0\]
rlabel metal2 48832 17752 48832 17752 0 spi.data_out_buff\[1\]
rlabel metal2 51016 14728 51016 14728 0 spi.data_out_buff\[2\]
rlabel metal2 52024 13944 52024 13944 0 spi.data_out_buff\[3\]
rlabel metal3 52304 19880 52304 19880 0 spi.data_out_buff\[4\]
rlabel metal2 50344 24248 50344 24248 0 spi.data_out_buff\[5\]
rlabel metal2 50344 26600 50344 26600 0 spi.data_out_buff\[6\]
rlabel metal2 48272 23688 48272 23688 0 spi.data_out_buff\[7\]
rlabel metal2 33824 9800 33824 9800 0 spi.div_counter\[0\]
rlabel metal2 34664 12880 34664 12880 0 spi.div_counter\[1\]
rlabel metal2 33712 15400 33712 15400 0 spi.div_counter\[2\]
rlabel metal2 39144 16828 39144 16828 0 spi.div_counter\[3\]
rlabel metal2 40936 13272 40936 13272 0 spi.div_counter\[4\]
rlabel metal2 36904 6216 36904 6216 0 spi.div_counter\[5\]
rlabel metal2 39592 16800 39592 16800 0 spi.div_counter\[6\]
rlabel metal2 39256 5824 39256 5824 0 spi.div_counter\[7\]
rlabel metal2 38696 21672 38696 21672 0 spi.divisor\[0\]
rlabel metal2 37352 22176 37352 22176 0 spi.divisor\[1\]
rlabel metal2 39368 16016 39368 16016 0 spi.divisor\[2\]
rlabel metal2 38696 18200 38696 18200 0 spi.divisor\[3\]
rlabel metal2 40264 16912 40264 16912 0 spi.divisor\[4\]
rlabel metal2 38808 28952 38808 28952 0 spi.divisor\[5\]
rlabel metal3 40488 23576 40488 23576 0 spi.divisor\[6\]
rlabel metal2 39760 35560 39760 35560 0 spi.divisor\[7\]
rlabel metal3 35504 21560 35504 21560 0 spi.dout\[0\]
rlabel metal2 31024 20552 31024 20552 0 spi.dout\[1\]
rlabel metal2 24248 13944 24248 13944 0 spi.dout\[2\]
rlabel metal2 28224 16744 28224 16744 0 spi.dout\[3\]
rlabel metal3 24416 17080 24416 17080 0 spi.dout\[4\]
rlabel metal2 23968 21784 23968 21784 0 spi.dout\[5\]
rlabel metal2 24024 20720 24024 20720 0 spi.dout\[6\]
rlabel metal2 27216 22456 27216 22456 0 spi.dout\[7\]
rlabel metal2 20328 19768 20328 19768 0 uart.busy
rlabel metal3 5320 13720 5320 13720 0 uart.counter\[0\]
rlabel metal2 5992 12880 5992 12880 0 uart.counter\[1\]
rlabel metal2 5208 11704 5208 11704 0 uart.counter\[2\]
rlabel metal2 5656 10416 5656 10416 0 uart.counter\[3\]
rlabel metal3 8400 7336 8400 7336 0 uart.data_buff\[0\]
rlabel metal2 10248 8372 10248 8372 0 uart.data_buff\[1\]
rlabel metal2 13160 7728 13160 7728 0 uart.data_buff\[2\]
rlabel metal2 14840 6384 14840 6384 0 uart.data_buff\[3\]
rlabel metal2 17528 8624 17528 8624 0 uart.data_buff\[4\]
rlabel metal2 19544 10192 19544 10192 0 uart.data_buff\[5\]
rlabel metal2 21672 15148 21672 15148 0 uart.data_buff\[6\]
rlabel metal2 20216 16912 20216 16912 0 uart.data_buff\[7\]
rlabel metal2 15568 18312 15568 18312 0 uart.data_buff\[8\]
rlabel metal2 12656 16184 12656 16184 0 uart.data_buff\[9\]
rlabel metal2 16296 29176 16296 29176 0 uart.div_counter\[0\]
rlabel metal3 16660 30184 16660 30184 0 uart.div_counter\[10\]
rlabel metal2 15960 32032 15960 32032 0 uart.div_counter\[11\]
rlabel metal3 16184 29288 16184 29288 0 uart.div_counter\[12\]
rlabel metal2 7560 22624 7560 22624 0 uart.div_counter\[13\]
rlabel metal2 18536 23632 18536 23632 0 uart.div_counter\[14\]
rlabel metal2 16408 21840 16408 21840 0 uart.div_counter\[15\]
rlabel metal2 19656 28784 19656 28784 0 uart.div_counter\[1\]
rlabel metal2 15624 26684 15624 26684 0 uart.div_counter\[2\]
rlabel metal2 16856 24416 16856 24416 0 uart.div_counter\[3\]
rlabel metal3 10528 34104 10528 34104 0 uart.div_counter\[4\]
rlabel metal2 12488 36400 12488 36400 0 uart.div_counter\[5\]
rlabel metal3 8176 35672 8176 35672 0 uart.div_counter\[6\]
rlabel metal3 10920 35896 10920 35896 0 uart.div_counter\[7\]
rlabel metal2 9464 25424 9464 25424 0 uart.div_counter\[8\]
rlabel metal2 8568 28224 8568 28224 0 uart.div_counter\[9\]
rlabel metal2 18312 26208 18312 26208 0 uart.divisor\[0\]
rlabel metal3 18928 37352 18928 37352 0 uart.divisor\[10\]
rlabel metal2 16296 34776 16296 34776 0 uart.divisor\[11\]
rlabel metal2 18312 33264 18312 33264 0 uart.divisor\[12\]
rlabel metal2 21896 32200 21896 32200 0 uart.divisor\[13\]
rlabel metal2 20160 24584 20160 24584 0 uart.divisor\[14\]
rlabel metal2 15568 36456 15568 36456 0 uart.divisor\[15\]
rlabel metal2 21112 37128 21112 37128 0 uart.divisor\[1\]
rlabel metal2 16968 30520 16968 30520 0 uart.divisor\[2\]
rlabel metal2 18816 28728 18816 28728 0 uart.divisor\[3\]
rlabel metal2 22008 34776 22008 34776 0 uart.divisor\[4\]
rlabel metal2 16744 36680 16744 36680 0 uart.divisor\[5\]
rlabel metal2 16072 35784 16072 35784 0 uart.divisor\[6\]
rlabel metal2 25368 35448 25368 35448 0 uart.divisor\[7\]
rlabel metal2 19096 25088 19096 25088 0 uart.divisor\[8\]
rlabel metal3 20104 35672 20104 35672 0 uart.divisor\[9\]
rlabel metal2 38808 39704 38808 39704 0 uart.dout\[0\]
rlabel metal3 33096 39368 33096 39368 0 uart.dout\[1\]
rlabel metal2 33152 41272 33152 41272 0 uart.dout\[2\]
rlabel metal2 41944 40320 41944 40320 0 uart.dout\[3\]
rlabel metal2 44632 41608 44632 41608 0 uart.dout\[4\]
rlabel metal2 44968 39256 44968 39256 0 uart.dout\[5\]
rlabel metal2 45136 38920 45136 38920 0 uart.dout\[6\]
rlabel metal2 40488 36792 40488 36792 0 uart.dout\[7\]
rlabel metal2 43512 20888 43512 20888 0 uart.has_byte
rlabel metal2 35056 42616 35056 42616 0 uart.receive_buff\[0\]
rlabel metal2 35336 50624 35336 50624 0 uart.receive_buff\[1\]
rlabel metal2 37016 50540 37016 50540 0 uart.receive_buff\[2\]
rlabel metal2 39816 49336 39816 49336 0 uart.receive_buff\[3\]
rlabel metal2 45584 49672 45584 49672 0 uart.receive_buff\[4\]
rlabel metal2 46312 46088 46312 46088 0 uart.receive_buff\[5\]
rlabel metal2 44240 44408 44240 44408 0 uart.receive_buff\[6\]
rlabel metal2 40376 46592 40376 46592 0 uart.receive_buff\[7\]
rlabel metal2 48832 49000 48832 49000 0 uart.receive_counter\[0\]
rlabel metal2 48888 46872 48888 46872 0 uart.receive_counter\[1\]
rlabel metal3 51128 49896 51128 49896 0 uart.receive_counter\[2\]
rlabel metal2 48888 45248 48888 45248 0 uart.receive_counter\[3\]
rlabel metal2 24248 41888 24248 41888 0 uart.receive_div_counter\[0\]
rlabel metal2 17864 43512 17864 43512 0 uart.receive_div_counter\[10\]
rlabel metal3 16128 46648 16128 46648 0 uart.receive_div_counter\[11\]
rlabel metal2 10528 44408 10528 44408 0 uart.receive_div_counter\[12\]
rlabel metal2 11592 45024 11592 45024 0 uart.receive_div_counter\[13\]
rlabel metal2 10920 40768 10920 40768 0 uart.receive_div_counter\[14\]
rlabel metal2 14728 39088 14728 39088 0 uart.receive_div_counter\[15\]
rlabel metal2 20328 40320 20328 40320 0 uart.receive_div_counter\[1\]
rlabel metal2 24584 39368 24584 39368 0 uart.receive_div_counter\[2\]
rlabel metal3 20776 40376 20776 40376 0 uart.receive_div_counter\[3\]
rlabel metal2 19712 50680 19712 50680 0 uart.receive_div_counter\[4\]
rlabel metal2 24808 46592 24808 46592 0 uart.receive_div_counter\[5\]
rlabel metal2 29176 50568 29176 50568 0 uart.receive_div_counter\[6\]
rlabel metal2 26096 48104 26096 48104 0 uart.receive_div_counter\[7\]
rlabel metal2 28504 42168 28504 42168 0 uart.receive_div_counter\[8\]
rlabel metal2 19432 45640 19432 45640 0 uart.receive_div_counter\[9\]
rlabel metal2 34216 44800 34216 44800 0 uart.receiving
rlabel metal3 45304 28840 45304 28840 0 uart_ien
rlabel metal2 13776 49000 13776 49000 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 55000 55000
<< end >>
