// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack_ptr[0] ;
 wire \as2650.stack_ptr[1] ;
 wire \as2650.stack_ptr[2] ;
 wire net90;
 wire clknet_leaf_0_wb_clk_i;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net91;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net92;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net93;
 wire net94;
 wire net79;
 wire net84;
 wire net80;
 wire net81;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net82;
 wire net83;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3588_ (.I(net53),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3589_ (.I(\as2650.ins_reg[1] ),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3590_ (.I(_3125_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3591_ (.I(_3126_),
    .Z(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3592_ (.I(_3127_),
    .Z(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3593_ (.I(\as2650.ins_reg[0] ),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3594_ (.I(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3595_ (.I(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3596_ (.I(_3131_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3597_ (.A1(_3128_),
    .A2(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3598_ (.I(_3133_),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3599_ (.A1(\as2650.halted ),
    .A2(net10),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3600_ (.I(\as2650.psl[4] ),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3601_ (.I(_3136_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3602_ (.I(_3137_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3603_ (.I(_3138_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3604_ (.I(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3605_ (.I(_3140_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3606_ (.I(\as2650.ins_reg[1] ),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3607_ (.I(_3142_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(\as2650.ins_reg[0] ),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3609_ (.A1(_3143_),
    .A2(_3144_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3610_ (.I(_3145_),
    .Z(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3611_ (.A1(_3141_),
    .A2(_3146_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3612_ (.A1(_3135_),
    .A2(_3147_),
    .Z(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3613_ (.I(_3148_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3614_ (.I(\as2650.cycle[0] ),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3615_ (.I(_3150_),
    .Z(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3616_ (.I(\as2650.cycle[1] ),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3617_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3618_ (.A1(\as2650.cycle[3] ),
    .A2(\as2650.cycle[2] ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3619_ (.A1(_3153_),
    .A2(_3154_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_3152_),
    .A2(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3621_ (.A1(_3151_),
    .A2(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3622_ (.I(_3157_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3623_ (.I(\as2650.ins_reg[3] ),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3624_ (.I(\as2650.ins_reg[2] ),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3625_ (.I(_3160_),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3626_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3627_ (.A1(\as2650.ins_reg[5] ),
    .A2(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3628_ (.I(_3163_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3629_ (.A1(_3161_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3630_ (.A1(_3159_),
    .A2(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3631_ (.A1(_3149_),
    .A2(_3158_),
    .A3(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3632_ (.I(_3167_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3633_ (.I(_3168_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3634_ (.I(_3135_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3635_ (.I(_3170_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3636_ (.I(_3147_),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3637_ (.I(_3155_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3638_ (.I(\as2650.cycle[1] ),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3639_ (.A1(_3174_),
    .A2(_3150_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3640_ (.A1(_3173_),
    .A2(_3175_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3641_ (.I(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3642_ (.I(_3177_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3643_ (.I(\as2650.ins_reg[3] ),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3644_ (.I(_3179_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3645_ (.I(_3180_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3646_ (.I(\as2650.ins_reg[2] ),
    .Z(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3647_ (.I(\as2650.ins_reg[4] ),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3648_ (.I(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(_3184_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3650_ (.I(\as2650.ins_reg[5] ),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3651_ (.I(_3186_),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(\as2650.ins_reg[6] ),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3653_ (.I(\as2650.ins_reg[7] ),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3654_ (.I(_3189_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3655_ (.A1(_3188_),
    .A2(_3190_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3656_ (.A1(_3182_),
    .A2(_3185_),
    .A3(_3187_),
    .A4(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3657_ (.A1(_3181_),
    .A2(_3192_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3658_ (.I(_3185_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3659_ (.I(\as2650.cycle[7] ),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3660_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3661_ (.I(_3152_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3662_ (.I(\as2650.cycle[0] ),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3663_ (.A1(_3197_),
    .A2(_3198_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3664_ (.A1(\as2650.cycle[6] ),
    .A2(_3154_),
    .A3(_3199_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3665_ (.A1(_3196_),
    .A2(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3666_ (.A1(_3195_),
    .A2(_3201_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3667_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3668_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3669_ (.A1(_3203_),
    .A2(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3670_ (.A1(_3194_),
    .A2(_3202_),
    .A3(_3205_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3671_ (.I(\as2650.ins_reg[3] ),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3672_ (.I(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3673_ (.I(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3674_ (.I(\as2650.ins_reg[4] ),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3675_ (.I(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3676_ (.I(_3211_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3677_ (.I(_3188_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3678_ (.I(_3157_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3679_ (.A1(_3209_),
    .A2(_3212_),
    .A3(_3213_),
    .A4(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3680_ (.A1(_3178_),
    .A2(_3193_),
    .B(_3206_),
    .C(_3215_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3681_ (.A1(_3172_),
    .A2(_3216_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(\as2650.ins_reg[7] ),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3683_ (.I(_3218_),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3684_ (.I(_3186_),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3685_ (.A1(_3161_),
    .A2(_3210_),
    .A3(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3686_ (.A1(_3219_),
    .A2(_3221_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3687_ (.I(_3222_),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3688_ (.I(_3153_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3689_ (.I(\as2650.cycle[3] ),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3690_ (.I(\as2650.cycle[2] ),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3691_ (.A1(_3152_),
    .A2(_3150_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3692_ (.A1(_3225_),
    .A2(_3226_),
    .A3(_3227_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3693_ (.A1(_3224_),
    .A2(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3694_ (.A1(_3209_),
    .A2(_3229_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3695_ (.A1(_3172_),
    .A2(_3223_),
    .A3(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3696_ (.I(_3211_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3697_ (.I(\as2650.addr_buff[5] ),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3698_ (.I(\as2650.addr_buff[6] ),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3699_ (.A1(_3233_),
    .A2(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3700_ (.I(_3235_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3701_ (.A1(_3232_),
    .A2(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3702_ (.I(_3237_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3703_ (.A1(\as2650.cycle[7] ),
    .A2(_3196_),
    .A3(_3200_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3704_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3239_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3705_ (.I(_3240_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3706_ (.A1(_3147_),
    .A2(_3238_),
    .A3(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3707_ (.A1(_3217_),
    .A2(_3231_),
    .A3(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3708_ (.A1(_3171_),
    .A2(_3243_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3709_ (.I(_3149_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3710_ (.I(_3158_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3711_ (.I(_3246_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3712_ (.I(\as2650.ins_reg[6] ),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3713_ (.I(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3714_ (.I(_3190_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3715_ (.A1(_3187_),
    .A2(_3249_),
    .A3(_3250_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3716_ (.I(_3210_),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3717_ (.A1(_3179_),
    .A2(_3160_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3718_ (.I(_3253_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3719_ (.I(_3254_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3720_ (.A1(_3252_),
    .A2(_3255_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3721_ (.A1(_3245_),
    .A2(_3247_),
    .A3(_3251_),
    .A4(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3722_ (.I(_3141_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3723_ (.I(_3252_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3724_ (.I(_3259_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3725_ (.I(\as2650.halted ),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3726_ (.I(net10),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3727_ (.A1(_3261_),
    .A2(_3262_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3728_ (.I(_3263_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3729_ (.A1(_3260_),
    .A2(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3730_ (.I(_3146_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3731_ (.I(_3205_),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3732_ (.A1(\as2650.ins_reg[3] ),
    .A2(\as2650.ins_reg[2] ),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3733_ (.I(_3268_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3734_ (.I(_3269_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3735_ (.I(_3270_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3736_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3737_ (.I(_3272_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3738_ (.I(\as2650.ins_reg[5] ),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3739_ (.A1(_3274_),
    .A2(_3248_),
    .A3(_3189_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3740_ (.A1(_3266_),
    .A2(_3267_),
    .A3(_3273_),
    .A4(_3275_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3741_ (.I(_3225_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3742_ (.A1(_3277_),
    .A2(_3226_),
    .A3(_3153_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3743_ (.A1(_3152_),
    .A2(_3150_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3744_ (.A1(_3278_),
    .A2(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3745_ (.I(_3280_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3746_ (.A1(_3265_),
    .A2(_3276_),
    .A3(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3747_ (.A1(_3258_),
    .A2(_3282_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3748_ (.A1(_3169_),
    .A2(_3244_),
    .A3(_3257_),
    .A4(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3749_ (.I(_3284_),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3750_ (.A1(_3134_),
    .A2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3751_ (.I(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3752_ (.I(\as2650.psl[4] ),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3753_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123_2[1][0] ),
    .S(_3288_),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3754_ (.A1(\as2650.r0[0] ),
    .A2(_3125_),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3755_ (.A1(_3126_),
    .A2(_3289_),
    .B(_3290_),
    .C(_3129_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _3756_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123[2][0] ),
    .I2(\as2650.r123_2[0][0] ),
    .I3(\as2650.r123_2[2][0] ),
    .S0(_3125_),
    .S1(_3288_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3757_ (.A1(\as2650.ins_reg[0] ),
    .A2(_3292_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3758_ (.A1(_3291_),
    .A2(_3293_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3759_ (.I(_3294_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3760_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3761_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3762_ (.A1(_3297_),
    .A2(_3204_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3763_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3764_ (.A1(_3203_),
    .A2(_3299_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3765_ (.A1(_3298_),
    .A2(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3766_ (.A1(_3296_),
    .A2(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3767_ (.I(_3302_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3768_ (.I(_3260_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3769_ (.I(_3195_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3770_ (.I(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3771_ (.I(_3201_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3772_ (.A1(_3306_),
    .A2(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3773_ (.A1(_3297_),
    .A2(_3299_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3774_ (.I(_3309_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3775_ (.A1(_3304_),
    .A2(_3308_),
    .A3(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3776_ (.A1(_3245_),
    .A2(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3777_ (.I(_3312_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3778_ (.I(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3779_ (.I(_3312_),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3780_ (.I(\as2650.r0[0] ),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3781_ (.I(_3316_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3782_ (.A1(_3251_),
    .A2(_3256_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3783_ (.A1(_3177_),
    .A2(_3318_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(_3149_),
    .A2(_3319_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3785_ (.I(_3320_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3786_ (.I(_3321_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3787_ (.I(_3167_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3788_ (.I(_3323_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3789_ (.I(\as2650.psl[3] ),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3790_ (.I(_3325_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3791_ (.A1(\as2650.r0[7] ),
    .A2(_3145_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3792_ (.I(_3137_),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3793_ (.I(_3328_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3794_ (.A1(_3139_),
    .A2(\as2650.r123[0][7] ),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3795_ (.I(_3125_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3796_ (.I(_3331_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3797_ (.A1(_3332_),
    .A2(_3132_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3798_ (.A1(_3329_),
    .A2(\as2650.r123_2[0][7] ),
    .B(_3330_),
    .C(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3799_ (.I(_3329_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3800_ (.I(\as2650.ins_reg[0] ),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3801_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3802_ (.A1(_3128_),
    .A2(_3337_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3803_ (.A1(_3139_),
    .A2(\as2650.r123[1][7] ),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3804_ (.A1(_3335_),
    .A2(\as2650.r123_2[1][7] ),
    .B(_3338_),
    .C(_3339_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3805_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_3139_),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3806_ (.A1(_3133_),
    .A2(_3341_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3807_ (.A1(_3327_),
    .A2(_3334_),
    .A3(_3340_),
    .A4(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3808_ (.I(_3343_),
    .Z(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3809_ (.I(_3344_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3810_ (.I(\as2650.carry ),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3811_ (.A1(\as2650.psl[3] ),
    .A2(_3346_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3812_ (.A1(_3326_),
    .A2(_3345_),
    .B(_3347_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3813_ (.A1(_3207_),
    .A2(_3176_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3814_ (.A1(_3192_),
    .A2(_3349_),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3815_ (.A1(_3149_),
    .A2(_3350_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3816_ (.I(_3351_),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3817_ (.I(_3352_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3818_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123_2[1][1] ),
    .S(_3288_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3819_ (.A1(\as2650.r0[1] ),
    .A2(_3331_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3820_ (.A1(_3126_),
    .A2(_3354_),
    .B(_3355_),
    .C(_3130_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3821_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123[2][1] ),
    .I2(\as2650.r123_2[0][1] ),
    .I3(\as2650.r123_2[2][1] ),
    .S0(_3142_),
    .S1(_3136_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3822_ (.A1(_3144_),
    .A2(_3357_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3823_ (.A1(_3356_),
    .A2(_3358_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3824_ (.I(_3359_),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3825_ (.I(_3360_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3826_ (.I(_3361_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3827_ (.A1(_3174_),
    .A2(_3198_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3828_ (.A1(_3173_),
    .A2(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3829_ (.A1(_3207_),
    .A2(_3364_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3830_ (.A1(_3148_),
    .A2(_3365_),
    .A3(_3222_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_3366_),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3832_ (.A1(_3291_),
    .A2(_3293_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3833_ (.I(_3368_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3834_ (.A1(_3162_),
    .A2(_3369_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3835_ (.I(net5),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3836_ (.I(_3371_),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3837_ (.I(_3372_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3838_ (.A1(_3373_),
    .A2(_3367_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3839_ (.A1(_3367_),
    .A2(_3370_),
    .B(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3840_ (.I(_3351_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3841_ (.A1(_3375_),
    .A2(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3842_ (.A1(_3353_),
    .A2(_3362_),
    .B(_3377_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3843_ (.A1(_3169_),
    .A2(_3378_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3844_ (.I(_3320_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3845_ (.A1(_3324_),
    .A2(_3348_),
    .B(_3379_),
    .C(_3380_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3846_ (.A1(_3170_),
    .A2(_3172_),
    .A3(_3238_),
    .A4(_3241_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3847_ (.I(_3382_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3848_ (.A1(_3317_),
    .A2(_3322_),
    .B(_3381_),
    .C(_3383_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3849_ (.I(\as2650.addr_buff[5] ),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3850_ (.A1(_3385_),
    .A2(\as2650.addr_buff[6] ),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3851_ (.I(\as2650.addr_buff[6] ),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3852_ (.A1(\as2650.addr_buff[5] ),
    .A2(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3853_ (.A1(_3386_),
    .A2(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3854_ (.A1(_3296_),
    .A2(_3389_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3855_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3856_ (.A1(_3170_),
    .A2(_3172_),
    .A3(_3238_),
    .A4(_3241_),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3857_ (.I(_3392_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3858_ (.A1(_3391_),
    .A2(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3859_ (.A1(_3315_),
    .A2(_3384_),
    .A3(_3394_),
    .ZN(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3860_ (.A1(_3303_),
    .A2(_3314_),
    .B(_3395_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3861_ (.I(_3250_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_3187_),
    .A2(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3863_ (.A1(_3213_),
    .A2(_3398_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3864_ (.I(_3399_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3865_ (.A1(_3220_),
    .A2(_3191_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3866_ (.I(_3401_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3867_ (.I(_3402_),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3868_ (.A1(_3316_),
    .A2(_3145_),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3869_ (.A1(_3332_),
    .A2(_3131_),
    .A3(_3289_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3870_ (.A1(_3336_),
    .A2(_3292_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3871_ (.I(\as2650.holding_reg[0] ),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3872_ (.A1(_3404_),
    .A2(_3405_),
    .A3(_3406_),
    .B(_3407_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3873_ (.A1(_3220_),
    .A2(_3249_),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3874_ (.I(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3875_ (.A1(_3407_),
    .A2(_3253_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3876_ (.I(\as2650.holding_reg[0] ),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _3877_ (.A1(_3291_),
    .A2(_3293_),
    .B(_3412_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3878_ (.A1(_3253_),
    .A2(_3295_),
    .B(_3411_),
    .C(_3413_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3879_ (.I(_3268_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3880_ (.I(_3294_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3881_ (.A1(_3407_),
    .A2(_3269_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3882_ (.A1(_3415_),
    .A2(_3416_),
    .B(_3417_),
    .C(_3413_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3883_ (.A1(_3414_),
    .A2(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3884_ (.A1(_3347_),
    .A2(_3419_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3885_ (.I(_3255_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3886_ (.I(_3368_),
    .Z(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3887_ (.I(_3422_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3888_ (.A1(_3412_),
    .A2(_3253_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3889_ (.A1(_3421_),
    .A2(_3423_),
    .B(_3424_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3890_ (.I(_3409_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3891_ (.A1(_3425_),
    .A2(_3426_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3892_ (.A1(_3186_),
    .A2(\as2650.ins_reg[6] ),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3893_ (.A1(_3218_),
    .A2(_3428_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3894_ (.I(_3429_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3895_ (.A1(_3410_),
    .A2(_3420_),
    .B(_3427_),
    .C(_3430_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3896_ (.I(\as2650.carry ),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3897_ (.A1(_3414_),
    .A2(_3418_),
    .B(\as2650.psl[3] ),
    .C(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3898_ (.A1(_3325_),
    .A2(_3432_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3899_ (.A1(_3434_),
    .A2(_3419_),
    .B(_3430_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3900_ (.I(_3191_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3901_ (.I(_3416_),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3902_ (.I(_3437_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3903_ (.A1(_3421_),
    .A2(_3438_),
    .B(_3411_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3904_ (.A1(_3274_),
    .A2(_3439_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3905_ (.A1(_3436_),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3906_ (.A1(_3433_),
    .A2(_3435_),
    .B(_3441_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3907_ (.A1(_3403_),
    .A2(_3408_),
    .B1(_3431_),
    .B2(_3442_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3908_ (.A1(_3419_),
    .A2(_3399_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3909_ (.A1(_3400_),
    .A2(_3443_),
    .B(_3444_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3910_ (.I(_3445_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3911_ (.A1(_3258_),
    .A2(_3282_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3912_ (.I0(_3396_),
    .I1(_3446_),
    .S(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3913_ (.I(net10),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3914_ (.A1(_3134_),
    .A2(_3284_),
    .B(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3915_ (.I(_3450_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3916_ (.A1(\as2650.r123[2][0] ),
    .A2(_3451_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3917_ (.A1(_3287_),
    .A2(_3448_),
    .B(_3452_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3918_ (.I(_3283_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3919_ (.A1(\as2650.holding_reg[1] ),
    .A2(_3269_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3920_ (.A1(_3269_),
    .A2(_3360_),
    .B(_3454_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3921_ (.A1(_3399_),
    .A2(_3455_),
    .ZN(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3922_ (.A1(_3356_),
    .A2(_3358_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3923_ (.I(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3924_ (.A1(\as2650.holding_reg[1] ),
    .A2(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3925_ (.I(\as2650.holding_reg[1] ),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3926_ (.A1(_3460_),
    .A2(_3458_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3927_ (.A1(_3459_),
    .A2(_3461_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3928_ (.A1(_3408_),
    .A2(_3433_),
    .B(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3929_ (.A1(_3459_),
    .A2(_3461_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3930_ (.A1(_3408_),
    .A2(_3433_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3931_ (.A1(_3218_),
    .A2(_3428_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3932_ (.A1(_3464_),
    .A2(_3465_),
    .B(_3466_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3933_ (.A1(_3254_),
    .A2(_3368_),
    .B(_3424_),
    .C(_3408_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3934_ (.A1(_3347_),
    .A2(_3468_),
    .B(_3414_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3935_ (.A1(_3464_),
    .A2(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3936_ (.A1(_3460_),
    .A2(_3255_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3937_ (.A1(_3255_),
    .A2(_3361_),
    .B(_3409_),
    .C(_3471_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3938_ (.A1(_3409_),
    .A2(_3470_),
    .B(_3472_),
    .C(_3429_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3939_ (.A1(_3463_),
    .A2(_3467_),
    .B(_3436_),
    .C(_3473_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3940_ (.I(_3457_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3941_ (.A1(_3460_),
    .A2(_3475_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3942_ (.A1(_3402_),
    .A2(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3943_ (.I(_3220_),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3944_ (.I(_3249_),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3945_ (.A1(_3479_),
    .A2(_3218_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3946_ (.A1(_3478_),
    .A2(_3480_),
    .A3(_3461_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3947_ (.A1(_3474_),
    .A2(_3477_),
    .A3(_3481_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3948_ (.I(_3482_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3949_ (.A1(_3456_),
    .A2(_3483_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3950_ (.I(_3283_),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3951_ (.A1(_3295_),
    .A2(_3359_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3952_ (.I(_3486_),
    .Z(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3953_ (.A1(_3385_),
    .A2(_3234_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3954_ (.A1(_3416_),
    .A2(_3386_),
    .B(_3488_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3955_ (.A1(_3487_),
    .A2(_3489_),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3956_ (.A1(_3487_),
    .A2(_3489_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3957_ (.A1(_3490_),
    .A2(_3491_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3958_ (.I(\as2650.r0[1] ),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3959_ (.I(_3493_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3960_ (.I(_3288_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3961_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123[2][2] ),
    .I2(\as2650.r123_2[0][2] ),
    .I3(\as2650.r123_2[2][2] ),
    .S0(_3142_),
    .S1(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3962_ (.A1(_3144_),
    .A2(_3496_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3963_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123_2[1][2] ),
    .S(_3136_),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3964_ (.A1(\as2650.r0[2] ),
    .A2(_3331_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3965_ (.A1(_3126_),
    .A2(_3498_),
    .B(_3499_),
    .C(_3130_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3966_ (.A1(_3497_),
    .A2(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3967_ (.I(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3968_ (.I(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3969_ (.I(_3503_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3970_ (.I(net6),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3971_ (.I(_3505_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3972_ (.I(_3506_),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3973_ (.A1(_3148_),
    .A2(_3365_),
    .A3(_3222_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3974_ (.I(_3508_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3975_ (.I(_3475_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3976_ (.A1(\as2650.ins_reg[4] ),
    .A2(_3275_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3977_ (.A1(_3296_),
    .A2(_3511_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3978_ (.A1(_3164_),
    .A2(_3437_),
    .B(_3512_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3979_ (.A1(_3510_),
    .A2(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_3509_),
    .A2(_3514_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3981_ (.A1(_3507_),
    .A2(_3509_),
    .B(_3376_),
    .C(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3982_ (.I(_3168_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3983_ (.A1(_3353_),
    .A2(_3504_),
    .B(_3516_),
    .C(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3984_ (.A1(_3324_),
    .A2(_3423_),
    .B(_3518_),
    .C(_3380_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3985_ (.A1(_3494_),
    .A2(_3322_),
    .B(_3382_),
    .C(_3519_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3986_ (.I(_3312_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3987_ (.A1(_3383_),
    .A2(_3492_),
    .B(_3520_),
    .C(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3988_ (.A1(_3297_),
    .A2(_3204_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3989_ (.A1(_3416_),
    .A2(_3298_),
    .B(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3990_ (.A1(_3487_),
    .A2(_3524_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3991_ (.A1(_3487_),
    .A2(_3524_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3992_ (.A1(_3525_),
    .A2(_3526_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3993_ (.A1(_3245_),
    .A2(_3311_),
    .A3(_3527_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3994_ (.A1(_3485_),
    .A2(_3522_),
    .A3(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3995_ (.A1(_3453_),
    .A2(_3484_),
    .B(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(\as2650.r123[2][1] ),
    .A2(_3451_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3997_ (.A1(_3287_),
    .A2(_3530_),
    .B(_3531_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3998_ (.A1(_3497_),
    .A2(_3500_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3999_ (.I(_3532_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4000_ (.I(_3533_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4001_ (.I(_3534_),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4002_ (.A1(_3423_),
    .A2(_3510_),
    .A3(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _4003_ (.A1(_3437_),
    .A2(_3361_),
    .B(_3503_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(_3203_),
    .A2(_3299_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4005_ (.A1(_3536_),
    .A2(_3537_),
    .B(_3538_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4006_ (.A1(_3422_),
    .A2(_3475_),
    .A3(_3533_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4007_ (.A1(_3437_),
    .A2(_3360_),
    .B(_3502_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4008_ (.A1(_3523_),
    .A2(_3540_),
    .A3(_3541_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4009_ (.I(_3301_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4010_ (.A1(_3543_),
    .A2(_3503_),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4011_ (.A1(_3539_),
    .A2(_3542_),
    .A3(_3544_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4012_ (.A1(\as2650.addr_buff[5] ),
    .A2(_3387_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4013_ (.A1(_3536_),
    .A2(_3537_),
    .B(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4014_ (.I(_3488_),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4015_ (.A1(_3548_),
    .A2(_3540_),
    .A3(_3541_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4016_ (.A1(_3546_),
    .A2(_3548_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4017_ (.A1(_3550_),
    .A2(_3535_),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4018_ (.A1(_3547_),
    .A2(_3549_),
    .A3(_3551_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4019_ (.A1(_3393_),
    .A2(_3552_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4020_ (.I(\as2650.r0[2] ),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4021_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123[2][3] ),
    .I2(\as2650.r123_2[0][3] ),
    .I3(\as2650.r123_2[2][3] ),
    .S0(_3142_),
    .S1(_3495_),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4022_ (.A1(_3144_),
    .A2(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4023_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123_2[1][3] ),
    .S(_3136_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4024_ (.A1(\as2650.r0[3] ),
    .A2(_3331_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4025_ (.A1(_3127_),
    .A2(_3557_),
    .B(_3558_),
    .C(_3130_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4026_ (.A1(_3556_),
    .A2(_3559_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4027_ (.I(_3560_),
    .Z(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4028_ (.I(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4029_ (.I(_3366_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4030_ (.I(_3458_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4031_ (.A1(_3163_),
    .A2(_3369_),
    .A3(_3564_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4032_ (.A1(_3369_),
    .A2(_3564_),
    .A3(_3511_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4033_ (.A1(_3503_),
    .A2(_3566_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4034_ (.I(net7),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4035_ (.I(_3568_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4036_ (.I(_3569_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4037_ (.A1(_3570_),
    .A2(_3563_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4038_ (.I(_3351_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4039_ (.A1(_3563_),
    .A2(_3567_),
    .B(_3571_),
    .C(_3572_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4040_ (.A1(_3353_),
    .A2(_3562_),
    .B(_3573_),
    .C(_3517_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4041_ (.A1(_3324_),
    .A2(_3362_),
    .B(_3574_),
    .C(_3380_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4042_ (.A1(_3554_),
    .A2(_3322_),
    .B(_3383_),
    .C(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4043_ (.A1(_3315_),
    .A2(_3553_),
    .A3(_3576_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4044_ (.A1(_3314_),
    .A2(_3545_),
    .B(_3577_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4045_ (.I(_3466_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4046_ (.I(\as2650.holding_reg[2] ),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4047_ (.A1(_3580_),
    .A2(_3533_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4048_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3533_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4049_ (.A1(_3581_),
    .A2(_3582_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4050_ (.I(_3583_),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4051_ (.A1(_3459_),
    .A2(_3463_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4052_ (.A1(_3584_),
    .A2(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4053_ (.A1(_3274_),
    .A2(_3213_),
    .A3(_3250_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4054_ (.I(_3587_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4055_ (.A1(_3455_),
    .A2(_3476_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4056_ (.A1(_3464_),
    .A2(_3469_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4057_ (.A1(_3584_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4058_ (.A1(_3415_),
    .A2(_3502_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4059_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3415_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4060_ (.A1(_3587_),
    .A2(_0266_),
    .B(_3430_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4061_ (.A1(_0261_),
    .A2(_0264_),
    .B(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4062_ (.A1(_3579_),
    .A2(_3586_),
    .B(_0268_),
    .C(_3480_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4063_ (.A1(_3478_),
    .A2(_3479_),
    .A3(_3397_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4064_ (.I(_3478_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4065_ (.A1(_3580_),
    .A2(_3535_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4066_ (.I(_3582_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4067_ (.A1(_0271_),
    .A2(_0272_),
    .B(_0273_),
    .C(_3480_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4068_ (.A1(_0270_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4069_ (.A1(_3399_),
    .A2(_3584_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4070_ (.A1(_0269_),
    .A2(_0275_),
    .B(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4071_ (.I(_0277_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4072_ (.I0(_3578_),
    .I1(_0278_),
    .S(_3447_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(\as2650.r123[2][2] ),
    .A2(_3451_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4074_ (.A1(_3287_),
    .A2(_0279_),
    .B(_0280_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4075_ (.I(_0270_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4076_ (.A1(_3556_),
    .A2(_3559_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4077_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4078_ (.I(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4079_ (.A1(_3584_),
    .A2(_0263_),
    .B1(_0266_),
    .B2(_0273_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4080_ (.A1(_0284_),
    .A2(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4081_ (.I(\as2650.holding_reg[3] ),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4082_ (.I(_0282_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4083_ (.I(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4084_ (.I(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4085_ (.A1(_3272_),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4086_ (.A1(_0287_),
    .A2(_3273_),
    .B(_3426_),
    .C(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4087_ (.I(_3430_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4088_ (.A1(_3410_),
    .A2(_0286_),
    .B(_0292_),
    .C(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4089_ (.A1(_3459_),
    .A2(_3463_),
    .A3(_0272_),
    .B(_0273_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4090_ (.A1(_0284_),
    .A2(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4091_ (.A1(_3579_),
    .A2(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(_3254_),
    .A2(_0288_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4093_ (.A1(\as2650.holding_reg[3] ),
    .A2(_3254_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4094_ (.A1(_0271_),
    .A2(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4095_ (.I(_3480_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4096_ (.A1(_0294_),
    .A2(_0297_),
    .B1(_0300_),
    .B2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4097_ (.A1(_0287_),
    .A2(_3561_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_3402_),
    .A2(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_0281_),
    .A2(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4100_ (.A1(_0281_),
    .A2(_0284_),
    .B1(_0302_),
    .B2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4101_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4102_ (.A1(_3540_),
    .A2(_0288_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4103_ (.A1(_3369_),
    .A2(_3564_),
    .A3(_3534_),
    .A4(_3561_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4104_ (.A1(_3296_),
    .A2(_3360_),
    .A3(_3502_),
    .B(_0288_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4105_ (.A1(_0309_),
    .A2(_0310_),
    .B(_3538_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4106_ (.A1(_3543_),
    .A2(_0290_),
    .B1(_0308_),
    .B2(_3300_),
    .C(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4107_ (.I(_0312_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4108_ (.I(_3321_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4109_ (.I(_3232_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4110_ (.I(\as2650.addr_buff[7] ),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4111_ (.I(\as2650.cycle[7] ),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4112_ (.A1(_0317_),
    .A2(_3307_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4113_ (.A1(_0315_),
    .A2(_0316_),
    .A3(_3236_),
    .A4(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4114_ (.A1(_3245_),
    .A2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4115_ (.I(_3535_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4116_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123_2[1][4] ),
    .S(_3137_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4117_ (.A1(\as2650.r0[4] ),
    .A2(_3332_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4118_ (.A1(_3127_),
    .A2(_0322_),
    .B(_0323_),
    .C(_3131_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4119_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123[2][4] ),
    .I2(\as2650.r123_2[0][4] ),
    .I3(\as2650.r123_2[2][4] ),
    .S0(_3143_),
    .S1(_3137_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(_3336_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4121_ (.A1(_0324_),
    .A2(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4122_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4123_ (.I(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4124_ (.I(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4125_ (.A1(_3163_),
    .A2(_3422_),
    .A3(_3564_),
    .A4(_3534_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4126_ (.A1(_3422_),
    .A2(_3475_),
    .A3(_3511_),
    .A4(_3534_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4127_ (.A1(_0331_),
    .A2(_0332_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4128_ (.A1(_0289_),
    .A2(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4129_ (.I(net8),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4130_ (.I(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4131_ (.I(_0336_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4132_ (.I(_0337_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4133_ (.A1(_0338_),
    .A2(_3366_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_3366_),
    .A2(_0334_),
    .B(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4135_ (.A1(_3352_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4136_ (.A1(_3376_),
    .A2(_0330_),
    .B(_0341_),
    .C(_3168_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4137_ (.A1(_3517_),
    .A2(_0321_),
    .B(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(_3257_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4139_ (.A1(\as2650.r0[3] ),
    .A2(_0314_),
    .B(_0320_),
    .C(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4140_ (.I(_3389_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4141_ (.A1(_0309_),
    .A2(_0310_),
    .B(_3546_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4142_ (.A1(_0346_),
    .A2(_0290_),
    .B1(_0308_),
    .B2(_3388_),
    .C(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4143_ (.I(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4144_ (.A1(_3392_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4145_ (.A1(_3313_),
    .A2(_0345_),
    .A3(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4146_ (.A1(_3521_),
    .A2(_0313_),
    .B(_0351_),
    .C(_3283_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4147_ (.I(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4148_ (.A1(_3447_),
    .A2(_0307_),
    .B(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4149_ (.A1(\as2650.r123[2][3] ),
    .A2(_3451_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4150_ (.A1(_3287_),
    .A2(_0354_),
    .B(_0355_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4151_ (.I(_3286_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4152_ (.A1(_3368_),
    .A2(_3458_),
    .A3(_3532_),
    .A4(_3560_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4153_ (.A1(_0357_),
    .A2(_0327_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4154_ (.A1(_3295_),
    .A2(_3359_),
    .A3(_3501_),
    .A4(_0282_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4155_ (.A1(_0359_),
    .A2(_0328_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4156_ (.A1(_3543_),
    .A2(_0328_),
    .B1(_0358_),
    .B2(_3300_),
    .C1(_3298_),
    .C2(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4157_ (.I(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4158_ (.I(\as2650.r0[4] ),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4159_ (.I(_0320_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4160_ (.I(_3562_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4161_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123[2][5] ),
    .I2(\as2650.r123_2[0][5] ),
    .I3(\as2650.r123_2[2][5] ),
    .S0(_3143_),
    .S1(_3495_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4162_ (.A1(_3336_),
    .A2(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4163_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123_2[1][5] ),
    .S(_3495_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4164_ (.A1(\as2650.r0[5] ),
    .A2(_3143_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4165_ (.A1(_3127_),
    .A2(_0368_),
    .B(_0369_),
    .C(_3131_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4166_ (.A1(_0367_),
    .A2(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4167_ (.I(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4168_ (.I(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4169_ (.I(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4170_ (.I(net9),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4171_ (.I(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4172_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4173_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4174_ (.A1(_3540_),
    .A2(_0289_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4175_ (.A1(_0331_),
    .A2(_0289_),
    .B1(_0379_),
    .B2(_3511_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4176_ (.A1(_0329_),
    .A2(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(_3508_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4178_ (.A1(_0378_),
    .A2(_3509_),
    .B(_3376_),
    .C(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4179_ (.A1(_3353_),
    .A2(_0374_),
    .B(_0383_),
    .C(_3323_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4180_ (.A1(_3324_),
    .A2(_0365_),
    .B(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(_3257_),
    .A2(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4182_ (.A1(_0363_),
    .A2(_3322_),
    .B(_0364_),
    .C(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4183_ (.A1(_3388_),
    .A2(_0358_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4184_ (.I(_3386_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4185_ (.A1(_0346_),
    .A2(_0329_),
    .B1(_0360_),
    .B2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4186_ (.A1(_0388_),
    .A2(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_3393_),
    .A2(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4188_ (.A1(_3521_),
    .A2(_0387_),
    .A3(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4189_ (.A1(_3314_),
    .A2(_0362_),
    .B(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4190_ (.I(_3400_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4191_ (.I(\as2650.holding_reg[4] ),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(_0324_),
    .A2(_0326_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4193_ (.A1(_0396_),
    .A2(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4194_ (.A1(_0396_),
    .A2(_0397_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4195_ (.A1(_0398_),
    .A2(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4196_ (.I(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4197_ (.I(_3403_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4198_ (.I(_3426_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4199_ (.A1(_3583_),
    .A2(_0284_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4200_ (.A1(\as2650.holding_reg[3] ),
    .A2(_3560_),
    .B(_0299_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4201_ (.A1(_0273_),
    .A2(_0266_),
    .A3(_0283_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4202_ (.A1(_0263_),
    .A2(_0404_),
    .B(_0405_),
    .C(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4203_ (.A1(_0401_),
    .A2(_0407_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4204_ (.I(_3421_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4205_ (.A1(_0396_),
    .A2(_3421_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4206_ (.A1(_0409_),
    .A2(_0330_),
    .B(_0410_),
    .C(_0403_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(_0293_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4208_ (.A1(_0403_),
    .A2(_0408_),
    .B(_0411_),
    .C(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4209_ (.A1(_0287_),
    .A2(_3562_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4210_ (.A1(_0414_),
    .A2(_0295_),
    .B(_0303_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4211_ (.A1(_0401_),
    .A2(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4212_ (.A1(\as2650.holding_reg[4] ),
    .A2(_3415_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4213_ (.A1(_3270_),
    .A2(_0327_),
    .B(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4214_ (.I(_0301_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4215_ (.A1(_3579_),
    .A2(_0416_),
    .B1(_0418_),
    .B2(_0419_),
    .C(_3403_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4216_ (.A1(_0402_),
    .A2(_0398_),
    .B1(_0413_),
    .B2(_0420_),
    .C(_3400_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4217_ (.A1(_0395_),
    .A2(_0401_),
    .B(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4218_ (.I(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4219_ (.I0(_0394_),
    .I1(_0423_),
    .S(_3447_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4220_ (.I(_3450_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4221_ (.A1(\as2650.r123[2][4] ),
    .A2(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4222_ (.A1(_0356_),
    .A2(_0424_),
    .B(_0426_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4223_ (.A1(_0367_),
    .A2(_0370_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4224_ (.I(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4225_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0428_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4226_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0428_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4227_ (.A1(_0429_),
    .A2(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4228_ (.I(_0430_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4229_ (.A1(_0429_),
    .A2(_0430_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4230_ (.A1(_0414_),
    .A2(_0295_),
    .B(_0398_),
    .C(_0303_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4231_ (.A1(_0399_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4232_ (.A1(_0433_),
    .A2(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4233_ (.A1(_0398_),
    .A2(_0418_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4234_ (.A1(_0400_),
    .A2(_0407_),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4235_ (.A1(_0431_),
    .A2(_0438_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4236_ (.I(\as2650.holding_reg[5] ),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4237_ (.A1(_3270_),
    .A2(_0371_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4238_ (.A1(_0440_),
    .A2(_3270_),
    .B(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4239_ (.A1(_3426_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4240_ (.A1(_3410_),
    .A2(_0439_),
    .B(_0443_),
    .C(_0293_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4241_ (.A1(_0271_),
    .A2(_0301_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4242_ (.A1(_0412_),
    .A2(_0436_),
    .B(_0444_),
    .C(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4243_ (.I(_3274_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4244_ (.I(_0428_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4245_ (.A1(_0440_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4246_ (.A1(_0447_),
    .A2(_0449_),
    .B(_0301_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4247_ (.A1(_3403_),
    .A2(_0432_),
    .B1(_0446_),
    .B2(_0450_),
    .C(_3400_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4248_ (.A1(_0395_),
    .A2(_0431_),
    .B(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4249_ (.I(_0452_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4250_ (.I(_3543_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4251_ (.A1(_0454_),
    .A2(_0373_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4252_ (.I(_3298_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4253_ (.I(_0397_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4254_ (.A1(_0359_),
    .A2(_0457_),
    .A3(_0428_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4255_ (.A1(_0309_),
    .A2(_0329_),
    .B(_0372_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4256_ (.A1(_0458_),
    .A2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4257_ (.A1(_0357_),
    .A2(_0328_),
    .B(_0371_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4258_ (.A1(_0397_),
    .A2(_0427_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4259_ (.A1(_0357_),
    .A2(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4260_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4261_ (.A1(_3523_),
    .A2(_0461_),
    .A3(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4262_ (.A1(_0456_),
    .A2(_0460_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4263_ (.A1(_0455_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4264_ (.A1(_3548_),
    .A2(_0461_),
    .A3(_0464_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4265_ (.A1(_0346_),
    .A2(_0372_),
    .B1(_0460_),
    .B2(_0389_),
    .C(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4266_ (.I(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4267_ (.I(\as2650.r0[5] ),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4268_ (.I(_0330_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4269_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_3138_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4270_ (.A1(_3133_),
    .A2(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4271_ (.A1(\as2650.r0[6] ),
    .A2(_3145_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4272_ (.A1(_3138_),
    .A2(\as2650.r123[0][6] ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4273_ (.A1(_3329_),
    .A2(\as2650.r123_2[0][6] ),
    .B(_3333_),
    .C(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4274_ (.A1(_3328_),
    .A2(\as2650.r123[1][6] ),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4275_ (.A1(_3329_),
    .A2(\as2650.r123_2[1][6] ),
    .B(_3338_),
    .C(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4276_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0477_),
    .A4(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4277_ (.I(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4278_ (.I(_0457_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4279_ (.A1(_0332_),
    .A2(_3561_),
    .A3(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4280_ (.A1(_3183_),
    .A2(_3275_),
    .A3(_0357_),
    .A4(_0462_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4281_ (.A1(_3164_),
    .A2(_0359_),
    .A3(_0457_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4282_ (.A1(_0483_),
    .A2(_0372_),
    .B(_0484_),
    .C(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4283_ (.A1(_3164_),
    .A2(_0359_),
    .A3(_0457_),
    .A4(_0448_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4284_ (.A1(_0486_),
    .A2(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(net1),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4286_ (.I(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4287_ (.A1(_0490_),
    .A2(_3367_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4288_ (.A1(_3563_),
    .A2(_0488_),
    .B(_0491_),
    .C(_3352_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4289_ (.A1(_3572_),
    .A2(_0481_),
    .B(_0492_),
    .C(_3323_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4290_ (.A1(_3169_),
    .A2(_0472_),
    .B(_0493_),
    .C(_3321_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4291_ (.A1(_0471_),
    .A2(_0314_),
    .B(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_0364_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4293_ (.A1(_3383_),
    .A2(_0470_),
    .B(_0496_),
    .C(_3521_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4294_ (.A1(_3314_),
    .A2(_0467_),
    .B(_0497_),
    .C(_3485_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4295_ (.A1(_3453_),
    .A2(_0453_),
    .B(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(\as2650.r123[2][5] ),
    .A2(_0425_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4297_ (.A1(_0356_),
    .A2(_0499_),
    .B(_0500_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(\as2650.holding_reg[6] ),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4299_ (.A1(_0501_),
    .A2(_0481_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4300_ (.I(_0480_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4301_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4302_ (.A1(_0502_),
    .A2(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4303_ (.I(_0505_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4304_ (.A1(_0399_),
    .A2(_0434_),
    .B(_0432_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4305_ (.A1(_0449_),
    .A2(_0506_),
    .A3(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4306_ (.A1(_0399_),
    .A2(_0429_),
    .A3(_0434_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4307_ (.A1(_0430_),
    .A2(_0506_),
    .A3(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4308_ (.A1(_0508_),
    .A2(_0510_),
    .B(_3579_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4309_ (.I(_3478_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4310_ (.A1(_0433_),
    .A2(_0437_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4311_ (.A1(_0429_),
    .A2(_0442_),
    .B(_0513_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4312_ (.A1(_0400_),
    .A2(_0407_),
    .A3(_0433_),
    .B(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4313_ (.A1(_0505_),
    .A2(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4314_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0477_),
    .A4(_0479_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4315_ (.A1(_3271_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4316_ (.A1(_0501_),
    .A2(_3271_),
    .B(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4317_ (.A1(_0261_),
    .A2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4318_ (.A1(_0261_),
    .A2(_0516_),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4319_ (.A1(_0512_),
    .A2(_0419_),
    .B1(_0412_),
    .B2(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4320_ (.A1(_0419_),
    .A2(_0504_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4321_ (.A1(_0511_),
    .A2(_0522_),
    .B(_0523_),
    .C(_0402_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4322_ (.A1(_0402_),
    .A2(_0502_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_0281_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4324_ (.A1(_0281_),
    .A2(_0506_),
    .B1(_0524_),
    .B2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4325_ (.I(_0527_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4326_ (.I(_0517_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4327_ (.I(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4328_ (.A1(_0458_),
    .A2(_0503_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4329_ (.A1(_0463_),
    .A2(_0503_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4330_ (.A1(_3523_),
    .A2(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4331_ (.A1(_0454_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_0456_),
    .C(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4332_ (.I(_0534_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(\as2650.r0[6] ),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4334_ (.A1(_0484_),
    .A2(_0487_),
    .A3(_0529_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4335_ (.I(net2),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4336_ (.I(_0538_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4337_ (.I(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4338_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4339_ (.A1(_0541_),
    .A2(_3367_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4340_ (.A1(_3563_),
    .A2(_0537_),
    .B(_0542_),
    .C(_3352_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4341_ (.A1(_3345_),
    .A2(_3572_),
    .B(_0543_),
    .C(_3323_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4342_ (.A1(_3169_),
    .A2(_0374_),
    .B(_0544_),
    .C(_3321_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4343_ (.A1(_0536_),
    .A2(_0314_),
    .B(_0364_),
    .C(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4344_ (.A1(_3548_),
    .A2(_0532_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4345_ (.A1(_0346_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_0389_),
    .C(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4346_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4347_ (.A1(_3393_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4348_ (.A1(_3313_),
    .A2(_0546_),
    .A3(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4349_ (.A1(_3315_),
    .A2(_0535_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4350_ (.A1(_3485_),
    .A2(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4351_ (.A1(_3453_),
    .A2(_0528_),
    .B(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4352_ (.A1(\as2650.r123[2][6] ),
    .A2(_0425_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4353_ (.A1(_0356_),
    .A2(_0554_),
    .B(_0555_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _4354_ (.A1(_3327_),
    .A2(_3334_),
    .A3(_3340_),
    .A4(_3342_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4355_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4357_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4358_ (.I(\as2650.holding_reg[7] ),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4359_ (.A1(_0560_),
    .A2(_3344_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4360_ (.A1(_0449_),
    .A2(_0505_),
    .A3(_0507_),
    .B(_0502_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4361_ (.A1(_0558_),
    .A2(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4362_ (.A1(_0504_),
    .A2(_0519_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4363_ (.A1(_0505_),
    .A2(_0515_),
    .B(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4364_ (.A1(_0557_),
    .A2(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4365_ (.I(_0556_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4366_ (.A1(_3272_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4367_ (.A1(\as2650.holding_reg[7] ),
    .A2(_3273_),
    .B(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_3410_),
    .A2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4369_ (.A1(_0403_),
    .A2(_0566_),
    .B(_0570_),
    .C(_0293_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4370_ (.A1(_0412_),
    .A2(_0563_),
    .B(_0571_),
    .C(_0445_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4371_ (.A1(\as2650.holding_reg[7] ),
    .A2(_3344_),
    .B(_0512_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(_0419_),
    .A2(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4373_ (.A1(_0402_),
    .A2(_0561_),
    .B1(_0572_),
    .B2(_0574_),
    .C(_0395_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4374_ (.A1(_0395_),
    .A2(_0559_),
    .B(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4375_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4376_ (.A1(_0458_),
    .A2(_0529_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4377_ (.A1(_0556_),
    .A2(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_0464_),
    .A2(_0529_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4379_ (.A1(_3343_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _4380_ (.A1(_0556_),
    .A2(_0454_),
    .B1(_0579_),
    .B2(_0456_),
    .C1(_0581_),
    .C2(_3300_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4381_ (.I(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(\as2650.r0[7] ),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4383_ (.I(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4384_ (.I(_0481_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4385_ (.A1(_3325_),
    .A2(_3423_),
    .B(_3347_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4386_ (.I(net3),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4387_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4388_ (.I0(_0484_),
    .I1(_0487_),
    .S(_0503_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4389_ (.A1(_3343_),
    .A2(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_3508_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4391_ (.A1(_0589_),
    .A2(_3509_),
    .B(_3351_),
    .C(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4392_ (.A1(_3572_),
    .A2(_0587_),
    .B(_0593_),
    .C(_3168_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4393_ (.A1(_3517_),
    .A2(_0586_),
    .B(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4394_ (.A1(_3380_),
    .A2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4395_ (.A1(_0585_),
    .A2(_0314_),
    .B(_0364_),
    .C(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4396_ (.A1(_3344_),
    .A2(_3550_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4397_ (.A1(_0389_),
    .A2(_0579_),
    .B1(_0581_),
    .B2(_3388_),
    .C(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4398_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4399_ (.A1(_3392_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4400_ (.A1(_3313_),
    .A2(_0597_),
    .A3(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4401_ (.A1(_3315_),
    .A2(_0583_),
    .B(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4402_ (.A1(_3485_),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4403_ (.A1(_3453_),
    .A2(_0577_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4404_ (.A1(\as2650.r123[2][7] ),
    .A2(_0425_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4405_ (.A1(_0356_),
    .A2(_0605_),
    .B(_0606_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(_3285_),
    .A2(_3338_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4407_ (.I(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4408_ (.A1(_3285_),
    .A2(_3338_),
    .B(_3449_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4410_ (.A1(\as2650.r123[1][0] ),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4411_ (.A1(_3448_),
    .A2(_0608_),
    .B(_0611_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4412_ (.A1(\as2650.r123[1][1] ),
    .A2(_0610_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4413_ (.A1(_3530_),
    .A2(_0608_),
    .B(_0612_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4414_ (.A1(\as2650.r123[1][2] ),
    .A2(_0610_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4415_ (.A1(_0279_),
    .A2(_0608_),
    .B(_0613_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4416_ (.A1(\as2650.r123[1][3] ),
    .A2(_0610_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4417_ (.A1(_0354_),
    .A2(_0608_),
    .B(_0614_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4418_ (.I(_0607_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4419_ (.I(_0609_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4420_ (.A1(\as2650.r123[1][4] ),
    .A2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4421_ (.A1(_0424_),
    .A2(_0615_),
    .B(_0617_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4422_ (.A1(\as2650.r123[1][5] ),
    .A2(_0616_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4423_ (.A1(_0499_),
    .A2(_0615_),
    .B(_0618_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4424_ (.A1(\as2650.r123[1][6] ),
    .A2(_0616_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4425_ (.A1(_0554_),
    .A2(_0615_),
    .B(_0619_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4426_ (.A1(\as2650.r123[1][7] ),
    .A2(_0616_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4427_ (.A1(_0605_),
    .A2(_0615_),
    .B(_0620_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4428_ (.I(_3197_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4429_ (.A1(_3277_),
    .A2(_3226_),
    .A3(_3224_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4430_ (.A1(_0621_),
    .A2(_3151_),
    .A3(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4431_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4432_ (.A1(_3141_),
    .A2(_3265_),
    .A3(_3276_),
    .A4(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4433_ (.I(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4434_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4435_ (.A1(_3335_),
    .A2(_3263_),
    .A3(_3146_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4436_ (.I(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4437_ (.A1(_3237_),
    .A2(_3240_),
    .A3(_0629_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4438_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4439_ (.I(_0631_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4440_ (.A1(_3319_),
    .A2(_0629_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4442_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_3214_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4444_ (.I(_3166_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4445_ (.I(_0629_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4446_ (.A1(_0636_),
    .A2(_0637_),
    .A3(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4447_ (.I(_3161_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4448_ (.A1(_0640_),
    .A2(_3252_),
    .A3(_3401_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4449_ (.A1(_3159_),
    .A2(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4450_ (.A1(_3158_),
    .A2(_0642_),
    .A3(_0628_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4451_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_3183_),
    .A2(_3186_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4453_ (.A1(_3182_),
    .A2(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4454_ (.A1(_3250_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_3128_),
    .A2(_3132_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4456_ (.A1(_3141_),
    .A2(_3170_),
    .A3(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4457_ (.A1(_3159_),
    .A2(_0647_),
    .A3(_3229_),
    .A4(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4459_ (.I(_0650_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4460_ (.A1(_3372_),
    .A2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4461_ (.A1(_3370_),
    .A2(_0651_),
    .B(_0643_),
    .C(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4462_ (.I(_3157_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4463_ (.A1(_0655_),
    .A2(_3166_),
    .A3(_0629_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4464_ (.I(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4465_ (.A1(_3510_),
    .A2(_0644_),
    .B(_0654_),
    .C(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4466_ (.A1(_3348_),
    .A2(_0639_),
    .B(_0658_),
    .C(_0634_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4467_ (.A1(_3317_),
    .A2(_0635_),
    .B(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4468_ (.A1(_0660_),
    .A2(_0631_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4469_ (.A1(_3311_),
    .A2(_0638_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4470_ (.A1(_3391_),
    .A2(_0632_),
    .B(_0661_),
    .C(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4471_ (.A1(_3206_),
    .A2(_0649_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(_3303_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4473_ (.A1(_0663_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4474_ (.I(_0625_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4475_ (.A1(_0666_),
    .A2(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4476_ (.A1(_3446_),
    .A2(_0627_),
    .B(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4477_ (.I(_3332_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4478_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4479_ (.I(_3337_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_0671_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4481_ (.A1(_0639_),
    .A2(_0625_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(_3209_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4483_ (.I(_3182_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4485_ (.I(_3364_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4486_ (.A1(_0677_),
    .A2(_3219_),
    .A3(_0678_),
    .A4(_0645_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4487_ (.A1(_0675_),
    .A2(_0679_),
    .A3(_0649_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4488_ (.A1(_0634_),
    .A2(_0680_),
    .A3(_0630_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4489_ (.A1(_3216_),
    .A2(_0638_),
    .B(_0674_),
    .C(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4490_ (.A1(_0673_),
    .A2(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4491_ (.I(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4492_ (.I0(_0669_),
    .I1(\as2650.r123_2[2][0] ),
    .S(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4493_ (.I(_0685_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4494_ (.I(_0684_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_0631_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4496_ (.I(_0662_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4497_ (.A1(_0319_),
    .A2(_0638_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_0634_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4499_ (.I(_0639_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4500_ (.I(_0643_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4501_ (.I(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(_0652_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(_3506_),
    .A2(_0651_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4504_ (.A1(_3514_),
    .A2(_0694_),
    .B(_0692_),
    .C(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4505_ (.A1(_0321_),
    .A2(_0693_),
    .B(_0696_),
    .C(_0657_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_0633_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4507_ (.A1(_3438_),
    .A2(_0691_),
    .B(_0697_),
    .C(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4508_ (.A1(_3493_),
    .A2(_0690_),
    .B(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4509_ (.A1(_0689_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4510_ (.A1(_3492_),
    .A2(_0687_),
    .B(_0688_),
    .C(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(_0664_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4512_ (.A1(_3527_),
    .A2(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4513_ (.A1(_0626_),
    .A2(_0702_),
    .A3(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4514_ (.A1(_3484_),
    .A2(_0627_),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(_0684_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4517_ (.A1(_0686_),
    .A2(_0706_),
    .B(_0708_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_0664_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4519_ (.I(_0698_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4520_ (.I(_3570_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4521_ (.I(_0650_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4522_ (.A1(_0711_),
    .A2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4523_ (.A1(_3567_),
    .A2(_0694_),
    .B(_0644_),
    .C(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_0656_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4525_ (.A1(_0365_),
    .A2(_0693_),
    .B(_0714_),
    .C(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4526_ (.A1(_3362_),
    .A2(_0691_),
    .B(_0716_),
    .C(_0635_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4527_ (.A1(_3554_),
    .A2(_0710_),
    .B(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_0631_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4529_ (.A1(_3552_),
    .A2(_0719_),
    .B(_0662_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4530_ (.A1(_0689_),
    .A2(_0718_),
    .B(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4531_ (.A1(_3545_),
    .A2(_0709_),
    .B(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4532_ (.I0(_0278_),
    .I1(_0722_),
    .S(_0667_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4533_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_0707_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4534_ (.A1(_0686_),
    .A2(_0723_),
    .B(_0724_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4535_ (.I(\as2650.r0[3] ),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(_3504_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_0657_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_0338_),
    .A2(_0652_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4539_ (.A1(_0334_),
    .A2(_0712_),
    .B(_0692_),
    .C(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4540_ (.A1(_0482_),
    .A2(_0644_),
    .B(_0729_),
    .C(_0657_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4541_ (.A1(_0726_),
    .A2(_0727_),
    .B(_0730_),
    .C(_0698_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4542_ (.A1(_0725_),
    .A2(_0690_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4543_ (.A1(_0689_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4544_ (.A1(_0349_),
    .A2(_0687_),
    .B(_0688_),
    .C(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4545_ (.A1(_0313_),
    .A2(_0703_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4546_ (.A1(_0626_),
    .A2(_0734_),
    .A3(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4547_ (.A1(_0307_),
    .A2(_0627_),
    .B(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_0683_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4549_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4550_ (.A1(_0686_),
    .A2(_0737_),
    .B(_0739_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4551_ (.A1(_0362_),
    .A2(_0709_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4552_ (.I(_0290_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4553_ (.A1(_0377_),
    .A2(_0651_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4554_ (.A1(_0381_),
    .A2(_0694_),
    .B(_0692_),
    .C(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4555_ (.A1(_0448_),
    .A2(_0693_),
    .B(_0743_),
    .C(_0715_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4556_ (.A1(_0741_),
    .A2(_0691_),
    .B(_0744_),
    .C(_0635_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4557_ (.A1(\as2650.r0[4] ),
    .A2(_0690_),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4558_ (.A1(_0632_),
    .A2(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4559_ (.A1(_0391_),
    .A2(_0687_),
    .B(_0688_),
    .C(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4560_ (.A1(_0667_),
    .A2(_0740_),
    .A3(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4561_ (.I(_0624_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4563_ (.A1(_3258_),
    .A2(_3265_),
    .A3(_3276_),
    .A4(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(_0423_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4565_ (.A1(_0749_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4566_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_0738_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4567_ (.A1(_0686_),
    .A2(_0754_),
    .B(_0755_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4568_ (.A1(_0467_),
    .A2(_0709_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4569_ (.I(_3177_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4570_ (.A1(_0757_),
    .A2(_3193_),
    .A3(_0649_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4571_ (.I(_0489_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4572_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4573_ (.I0(_0488_),
    .I1(_0760_),
    .S(_0712_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4574_ (.A1(_0481_),
    .A2(_0758_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4575_ (.A1(_0758_),
    .A2(_0761_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_0727_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4577_ (.A1(_0472_),
    .A2(_0727_),
    .B(_0764_),
    .C(_0710_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4578_ (.A1(_0471_),
    .A2(_0710_),
    .B(_0632_),
    .C(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4579_ (.I(_0719_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4580_ (.A1(_0470_),
    .A2(_0767_),
    .B(_0703_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4581_ (.A1(_0766_),
    .A2(_0768_),
    .B(_0752_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4582_ (.A1(_0453_),
    .A2(_0752_),
    .B1(_0756_),
    .B2(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4583_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_0738_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4584_ (.A1(_0707_),
    .A2(_0770_),
    .B(_0771_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4585_ (.I(_0374_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4586_ (.I(_3345_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(_0541_),
    .A2(_0712_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4588_ (.A1(_0537_),
    .A2(_0694_),
    .B(_0644_),
    .C(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4589_ (.A1(_0773_),
    .A2(_0693_),
    .B(_0775_),
    .C(_0715_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4590_ (.A1(_0772_),
    .A2(_0727_),
    .B(_0776_),
    .C(_0635_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4591_ (.A1(_0536_),
    .A2(_0710_),
    .B(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4592_ (.A1(_0549_),
    .A2(_0719_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4593_ (.A1(_0632_),
    .A2(_0778_),
    .B(_0779_),
    .C(_0664_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4594_ (.A1(_0535_),
    .A2(_0709_),
    .B(_0752_),
    .C(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4595_ (.A1(_0528_),
    .A2(_0667_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4596_ (.A1(_0781_),
    .A2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4597_ (.I0(_0783_),
    .I1(\as2650.r123_2[2][6] ),
    .S(_0684_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4598_ (.I(_0784_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4599_ (.I(_0530_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4600_ (.A1(_0591_),
    .A2(_0652_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4601_ (.A1(_0589_),
    .A2(_0651_),
    .B(_0758_),
    .C(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4602_ (.A1(_0587_),
    .A2(_0758_),
    .B(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(_0715_),
    .A2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4604_ (.A1(_0785_),
    .A2(_0691_),
    .B(_0789_),
    .C(_0698_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4605_ (.A1(_0585_),
    .A2(_0690_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_0719_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4607_ (.A1(_0600_),
    .A2(_0687_),
    .B(_0688_),
    .C(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4608_ (.A1(_0583_),
    .A2(_0703_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4609_ (.A1(_0626_),
    .A2(_0793_),
    .A3(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4610_ (.A1(_0577_),
    .A2(_0627_),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_0738_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4612_ (.A1(_0707_),
    .A2(_0796_),
    .B(_0797_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4613_ (.I(_3333_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_3180_),
    .A2(_3182_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4615_ (.I(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4616_ (.A1(_3436_),
    .A2(_0645_),
    .A3(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4617_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_0798_),
    .A2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4619_ (.I(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4620_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4621_ (.I(_3192_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4622_ (.A1(_0676_),
    .A2(_0271_),
    .A3(_3162_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4623_ (.A1(_0806_),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4624_ (.A1(_3221_),
    .A2(_0808_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4625_ (.I(_0640_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4626_ (.A1(_3183_),
    .A2(_3249_),
    .A3(_3190_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4627_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4628_ (.A1(_0810_),
    .A2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4629_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4630_ (.A1(_0673_),
    .A2(_0802_),
    .B(_0809_),
    .C(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4631_ (.I(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4632_ (.I(_0678_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4635_ (.A1(_0805_),
    .A2(_0816_),
    .B(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4636_ (.I(_3178_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4637_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4638_ (.I(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4639_ (.I(_0813_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4640_ (.I(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_3128_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4642_ (.A1(_3252_),
    .A2(_3271_),
    .A3(_3466_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4643_ (.A1(_0826_),
    .A2(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4644_ (.I(_0828_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4645_ (.A1(_0672_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4646_ (.I(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4647_ (.I(_0677_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4648_ (.I(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4649_ (.A1(_3187_),
    .A2(_0812_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4650_ (.I(_3174_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4651_ (.A1(_3224_),
    .A2(_3154_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4652_ (.I(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4653_ (.A1(_0835_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4654_ (.I(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_3261_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4656_ (.A1(_0833_),
    .A2(_0834_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4657_ (.A1(_0823_),
    .A2(_0825_),
    .A3(_0831_),
    .B(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4658_ (.A1(_0671_),
    .A2(_0827_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_3337_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4660_ (.A1(_0670_),
    .A2(_3272_),
    .A3(_0834_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4661_ (.A1(_0844_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4662_ (.I(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4663_ (.I(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4664_ (.A1(_0843_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4665_ (.A1(_3181_),
    .A2(_3211_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4666_ (.A1(_0621_),
    .A2(_0837_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4667_ (.A1(_0850_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_0821_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4669_ (.I(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4670_ (.I(_0824_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4671_ (.A1(_0854_),
    .A2(_0855_),
    .B(_0809_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4672_ (.I(_0677_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4673_ (.A1(\as2650.psl[6] ),
    .A2(_3337_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4674_ (.A1(\as2650.psl[7] ),
    .A2(_0670_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4675_ (.A1(_0858_),
    .A2(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4676_ (.A1(_3134_),
    .A2(_0812_),
    .A3(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(_0857_),
    .A2(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4679_ (.A1(_0849_),
    .A2(_0852_),
    .A3(_0856_),
    .A4(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4680_ (.A1(_0820_),
    .A2(_0842_),
    .A3(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4681_ (.A1(_3161_),
    .A2(_0811_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4682_ (.I(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4683_ (.I(_0636_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4684_ (.I(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4685_ (.A1(\as2650.r0[5] ),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4686_ (.I(_0490_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4687_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4689_ (.I(_0853_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4690_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_3266_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4692_ (.I(_0802_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4693_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4694_ (.A1(_0873_),
    .A2(_0876_),
    .A3(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4695_ (.A1(\as2650.psu[5] ),
    .A2(_0873_),
    .B(_0875_),
    .C(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4696_ (.A1(_0870_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4697_ (.A1(_0867_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4698_ (.I(_3262_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4699_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4700_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4701_ (.A1(\as2650.psu[5] ),
    .A2(_0865_),
    .B(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4702_ (.A1(_0865_),
    .A2(_0882_),
    .B(_0886_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4703_ (.I(\as2650.pc[0] ),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4704_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4705_ (.I(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4706_ (.I(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4707_ (.I(_0890_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(\as2650.stack_ptr[2] ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4710_ (.I(_0893_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4711_ (.I(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(\as2650.stack_ptr[1] ),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4713_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4714_ (.I(_0897_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4715_ (.I(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4716_ (.I(_0678_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4717_ (.A1(_3174_),
    .A2(_3278_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4718_ (.A1(_3151_),
    .A2(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4719_ (.I(_3198_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4720_ (.I(\as2650.cycle[2] ),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4721_ (.A1(_3225_),
    .A2(_0904_),
    .A3(_3224_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4722_ (.A1(_3197_),
    .A2(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4723_ (.A1(_0903_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4724_ (.A1(_0902_),
    .A2(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4725_ (.I(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4726_ (.A1(_0316_),
    .A2(_0623_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4727_ (.A1(_0909_),
    .A2(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4728_ (.A1(_0857_),
    .A2(_0900_),
    .B(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4729_ (.I(_3185_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4730_ (.I(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4731_ (.A1(_3398_),
    .A2(_0403_),
    .B(_0914_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4732_ (.A1(_3184_),
    .A2(_3188_),
    .A3(_3190_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4733_ (.A1(_3133_),
    .A2(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4734_ (.I(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4735_ (.A1(_3181_),
    .A2(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4736_ (.A1(_0912_),
    .A2(_0915_),
    .A3(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4737_ (.I(_3281_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_3207_),
    .A2(_0918_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4739_ (.A1(_0640_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4740_ (.I(_0923_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4741_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4742_ (.A1(_0512_),
    .A2(_0921_),
    .A3(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4743_ (.I(\as2650.stack_ptr[0] ),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4744_ (.I(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4745_ (.I(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4746_ (.A1(_0920_),
    .A2(_0926_),
    .B(_0929_),
    .C(_3264_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4747_ (.A1(_0895_),
    .A2(_0899_),
    .A3(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4748_ (.I(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4749_ (.I(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_0931_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4751_ (.A1(\as2650.stack[6][0] ),
    .A2(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4752_ (.A1(_0892_),
    .A2(_0933_),
    .B(_0935_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4753_ (.I(\as2650.pc[1] ),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4754_ (.I(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4756_ (.I(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(\as2650.stack[6][1] ),
    .A2(_0934_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4758_ (.A1(_0939_),
    .A2(_0933_),
    .B(_0940_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4759_ (.I(\as2650.pc[2] ),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4760_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4761_ (.I(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4762_ (.I(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4763_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4764_ (.A1(\as2650.stack[6][2] ),
    .A2(_0934_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4765_ (.A1(_0945_),
    .A2(_0933_),
    .B(_0946_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4766_ (.I(\as2650.pc[3] ),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4767_ (.I(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4768_ (.I(_0948_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4769_ (.I(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(\as2650.stack[6][3] ),
    .A2(_0934_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4772_ (.A1(_0951_),
    .A2(_0933_),
    .B(_0952_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4773_ (.I(\as2650.pc[4] ),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4774_ (.I(_0953_),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4775_ (.I(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4776_ (.I(_0932_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4777_ (.I(_0931_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(\as2650.stack[6][4] ),
    .A2(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4779_ (.A1(_0955_),
    .A2(_0956_),
    .B(_0958_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4780_ (.I(\as2650.pc[5] ),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4781_ (.I(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4782_ (.I(_0960_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4783_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4784_ (.A1(\as2650.stack[6][5] ),
    .A2(_0957_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4785_ (.A1(_0962_),
    .A2(_0956_),
    .B(_0963_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4786_ (.I(\as2650.pc[6] ),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4787_ (.I(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_0966_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(\as2650.stack[6][6] ),
    .A2(_0957_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4791_ (.A1(_0967_),
    .A2(_0956_),
    .B(_0968_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4792_ (.I(\as2650.pc[7] ),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4793_ (.I(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4795_ (.I(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4796_ (.A1(\as2650.stack[6][7] ),
    .A2(_0957_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4797_ (.A1(_0972_),
    .A2(_0956_),
    .B(_0973_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4798_ (.I(\as2650.pc[8] ),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4799_ (.I(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4800_ (.I(_0975_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4802_ (.I0(_0977_),
    .I1(\as2650.stack[6][8] ),
    .S(_0932_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4803_ (.I(_0978_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4804_ (.I(\as2650.pc[9] ),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4805_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4806_ (.I(_0980_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4807_ (.I(_0932_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_0931_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4809_ (.A1(\as2650.stack[6][9] ),
    .A2(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4810_ (.A1(_0981_),
    .A2(_0982_),
    .B(_0984_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4811_ (.I(\as2650.pc[10] ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4812_ (.I(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4813_ (.I(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4814_ (.A1(\as2650.stack[6][10] ),
    .A2(_0983_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4815_ (.A1(_0987_),
    .A2(_0982_),
    .B(_0988_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4816_ (.I(\as2650.pc[11] ),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4817_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(\as2650.stack[6][11] ),
    .A2(_0983_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4820_ (.A1(_0991_),
    .A2(_0982_),
    .B(_0992_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4821_ (.I(\as2650.pc[12] ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4823_ (.I(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4824_ (.A1(\as2650.stack[6][12] ),
    .A2(_0983_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4825_ (.A1(_0995_),
    .A2(_0982_),
    .B(_0996_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4826_ (.I(\as2650.psl[6] ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4827_ (.A1(_3178_),
    .A2(_0850_),
    .A3(_0813_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4828_ (.A1(_0836_),
    .A2(_3227_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4829_ (.I(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4830_ (.A1(_3436_),
    .A2(_0645_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4831_ (.A1(_0844_),
    .A2(_0800_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4832_ (.A1(_1000_),
    .A2(_1001_),
    .A3(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4833_ (.A1(_3194_),
    .A2(_0757_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4834_ (.I(_0622_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4835_ (.A1(_0835_),
    .A2(_0903_),
    .A3(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4836_ (.A1(_3364_),
    .A2(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4837_ (.A1(_1004_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4838_ (.A1(_0830_),
    .A2(_0998_),
    .B(_1003_),
    .C(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4839_ (.A1(_3180_),
    .A2(_0866_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4840_ (.A1(_3194_),
    .A2(_3158_),
    .A3(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4841_ (.A1(_3178_),
    .A2(_0642_),
    .B1(_0807_),
    .B2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4842_ (.A1(_0812_),
    .A2(_0800_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4843_ (.A1(_3259_),
    .A2(_3364_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4844_ (.A1(_1013_),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4845_ (.A1(_3266_),
    .A2(_3319_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4846_ (.A1(_3232_),
    .A2(_3177_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4847_ (.A1(_3219_),
    .A2(_0646_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4848_ (.A1(_3159_),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4849_ (.A1(_0409_),
    .A2(_1017_),
    .B(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4850_ (.A1(_1012_),
    .A2(_1015_),
    .A3(_1016_),
    .A4(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4851_ (.I(_3273_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4852_ (.A1(_0914_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4853_ (.A1(_0648_),
    .A2(_3318_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4854_ (.I(_3213_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4855_ (.I(_3219_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4856_ (.A1(_3212_),
    .A2(_0512_),
    .A3(_1025_),
    .A4(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4857_ (.A1(_3146_),
    .A2(_3402_),
    .A3(_3256_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_3157_),
    .A2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4859_ (.A1(_1023_),
    .A2(_1024_),
    .A3(_1027_),
    .A4(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4860_ (.A1(_3318_),
    .A2(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4861_ (.I(_3173_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4862_ (.A1(_0835_),
    .A2(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4863_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4865_ (.I(\as2650.halted ),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4866_ (.A1(_0757_),
    .A2(_1028_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4867_ (.A1(_1036_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4868_ (.A1(_1035_),
    .A2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_3156_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4870_ (.I(_0647_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4871_ (.A1(_3208_),
    .A2(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4872_ (.I(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4873_ (.A1(_1040_),
    .A2(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(_3208_),
    .A2(_3259_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4875_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4876_ (.A1(_1042_),
    .A2(_0843_),
    .B(_0636_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4877_ (.I(_3304_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4878_ (.A1(_1048_),
    .A2(_0447_),
    .A3(_3365_),
    .A4(_0815_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4879_ (.A1(_1044_),
    .A2(_1046_),
    .A3(_1047_),
    .A4(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4880_ (.I(_0999_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4881_ (.I(_1051_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4882_ (.A1(_0641_),
    .A2(_3165_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4883_ (.A1(_0646_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4884_ (.A1(_1054_),
    .A2(_1011_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4885_ (.A1(_0670_),
    .A2(_0827_),
    .B(_0845_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4886_ (.I(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4887_ (.A1(_1054_),
    .A2(_1057_),
    .A3(_0998_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4888_ (.I(_0829_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4889_ (.A1(_1052_),
    .A2(_1055_),
    .B1(_1058_),
    .B2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4890_ (.A1(_1039_),
    .A2(_1050_),
    .A3(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4891_ (.A1(_1009_),
    .A2(_1021_),
    .A3(_1031_),
    .A4(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4892_ (.I(_3275_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4893_ (.I(\as2650.psl[1] ),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4894_ (.A1(_0506_),
    .A2(_0558_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4895_ (.A1(_0401_),
    .A2(_0433_),
    .A3(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4896_ (.A1(_3418_),
    .A2(_3464_),
    .B(_0262_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4897_ (.A1(_0404_),
    .A2(_1067_),
    .B(_0405_),
    .C(_0406_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4898_ (.A1(_1066_),
    .A2(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4899_ (.A1(_0560_),
    .A2(_3345_),
    .B(_0569_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4900_ (.A1(_1069_),
    .A2(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4901_ (.A1(_1064_),
    .A2(_0559_),
    .A3(_1071_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4902_ (.A1(_0514_),
    .A2(_1065_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4903_ (.A1(_1064_),
    .A2(_0558_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4904_ (.A1(_0559_),
    .A2(_0564_),
    .B(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4905_ (.A1(_1073_),
    .A2(_1071_),
    .A3(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4906_ (.A1(_1063_),
    .A2(_1072_),
    .A3(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4907_ (.A1(_3419_),
    .A2(_3462_),
    .A3(_0404_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4908_ (.A1(_1066_),
    .A2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4909_ (.I(_3259_),
    .Z(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4910_ (.I(_1080_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4911_ (.A1(_1081_),
    .A2(_0868_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4912_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4913_ (.I(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4914_ (.I(_0576_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4915_ (.A1(_3456_),
    .A2(_3482_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4916_ (.A1(_3446_),
    .A2(_1086_),
    .A3(_0278_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4917_ (.A1(_0307_),
    .A2(_1087_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4918_ (.A1(_0422_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4919_ (.A1(_0452_),
    .A2(_0527_),
    .A3(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4920_ (.A1(_1063_),
    .A2(_1085_),
    .A3(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4921_ (.A1(_1077_),
    .A2(_1079_),
    .B(_1084_),
    .C(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4922_ (.I(_1081_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4923_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4924_ (.I(_0641_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_1095_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_3165_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4928_ (.I(_0845_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4929_ (.A1(_3554_),
    .A2(_3493_),
    .A3(_3316_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4930_ (.A1(\as2650.r0[6] ),
    .A2(\as2650.r0[5] ),
    .A3(\as2650.r0[4] ),
    .A4(\as2650.r0[3] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4931_ (.A1(_1100_),
    .A2(_1101_),
    .B(_0584_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4932_ (.I(_0536_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4933_ (.A1(_1103_),
    .A2(_1099_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4934_ (.I(_0636_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4935_ (.A1(_1099_),
    .A2(_1102_),
    .B(_1104_),
    .C(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4936_ (.I(_0757_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4937_ (.I(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4938_ (.I(_0541_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4939_ (.A1(\as2650.psl[6] ),
    .A2(_0541_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4940_ (.A1(_0826_),
    .A2(_1109_),
    .B(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4941_ (.A1(_0672_),
    .A2(_1108_),
    .A3(_0877_),
    .A4(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4942_ (.A1(_1098_),
    .A2(_1106_),
    .A3(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_0807_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4944_ (.A1(_1114_),
    .A2(_0586_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4945_ (.A1(_1114_),
    .A2(_3348_),
    .A3(_0464_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4946_ (.A1(_1113_),
    .A2(_1115_),
    .A3(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_3510_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4948_ (.A1(_0773_),
    .A2(_1118_),
    .A3(_0321_),
    .A4(_3562_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4949_ (.A1(_0462_),
    .A2(_0785_),
    .A3(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4950_ (.I(_1095_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4951_ (.A1(_0587_),
    .A2(_1120_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4952_ (.I(_3223_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4953_ (.A1(_1096_),
    .A2(_1117_),
    .B(_1122_),
    .C(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4954_ (.I(_0378_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4955_ (.I(_1109_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4956_ (.A1(_1125_),
    .A2(_0871_),
    .A3(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4957_ (.I(_3373_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_3507_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4959_ (.I(_0711_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4960_ (.I(_0338_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4961_ (.I(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4962_ (.A1(_1128_),
    .A2(_1129_),
    .A3(_1130_),
    .A4(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4963_ (.I(net3),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4964_ (.I(_1134_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4965_ (.I(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4966_ (.I(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4967_ (.I(_1041_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4968_ (.A1(_1127_),
    .A2(_1133_),
    .B(_1137_),
    .C(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4969_ (.A1(_1124_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4970_ (.I(_0567_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4971_ (.A1(_1141_),
    .A2(_0580_),
    .A3(_1027_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4972_ (.I(_0914_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4973_ (.A1(_1143_),
    .A2(_3397_),
    .A3(_3428_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4974_ (.A1(_0914_),
    .A2(_3247_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4975_ (.A1(_1144_),
    .A2(_1102_),
    .B(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4976_ (.A1(_1094_),
    .A2(_1140_),
    .B1(_1142_),
    .B2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4977_ (.A1(_1092_),
    .A2(_1147_),
    .B(_1062_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4978_ (.I(net10),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4979_ (.I(_1149_),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4980_ (.A1(_0997_),
    .A2(_1062_),
    .B(_1148_),
    .C(_1150_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4981_ (.I(_0884_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4982_ (.A1(_1063_),
    .A2(_1085_),
    .B(_1077_),
    .C(_0854_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4983_ (.A1(_0584_),
    .A2(_1093_),
    .A3(_1027_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4984_ (.I(_1004_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4985_ (.A1(_0773_),
    .A2(_1144_),
    .B(_1153_),
    .C(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4986_ (.I(_0589_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_1156_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4988_ (.I(_1041_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4989_ (.I(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(\as2650.psl[7] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4991_ (.I(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4992_ (.A1(_3569_),
    .A2(_3504_),
    .B1(_0741_),
    .B2(_0337_),
    .C1(_0373_),
    .C2(_0490_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4993_ (.A1(_0588_),
    .A2(_0567_),
    .B1(_3361_),
    .B2(_3506_),
    .C1(_0330_),
    .C2(_0377_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_0539_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4995_ (.I(_3132_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4996_ (.A1(_3211_),
    .A2(_3587_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4997_ (.A1(_1165_),
    .A2(_0799_),
    .A3(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4998_ (.A1(_3372_),
    .A2(_3438_),
    .B1(_0530_),
    .B2(_1164_),
    .C(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4999_ (.A1(_1162_),
    .A2(_1163_),
    .A3(_1168_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5000_ (.I(\as2650.overflow ),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5001_ (.I(_3505_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5002_ (.I(_1171_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5003_ (.I(_1172_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5004_ (.I(_0336_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5005_ (.I(_3372_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _5006_ (.A1(\as2650.psl[1] ),
    .A2(_1173_),
    .B1(_1174_),
    .B2(_3325_),
    .C1(_3432_),
    .C2(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5007_ (.A1(_1170_),
    .A2(_3569_),
    .B1(_0376_),
    .B2(_3335_),
    .C(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5008_ (.I(\as2650.psl[5] ),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5009_ (.A1(_1161_),
    .A2(_1134_),
    .B1(_0540_),
    .B2(_0997_),
    .C1(_0490_),
    .C2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5010_ (.A1(_1167_),
    .A2(_1177_),
    .A3(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5011_ (.A1(_0844_),
    .A2(_0800_),
    .A3(_1166_),
    .B(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5012_ (.I(\as2650.psu[7] ),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5013_ (.I(\as2650.psu[2] ),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5014_ (.I(_0375_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(net2),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5016_ (.I(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_1186_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5018_ (.A1(\as2650.psu[4] ),
    .A2(_1184_),
    .B1(_1187_),
    .B2(net27),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5019_ (.A1(\as2650.psu[1] ),
    .A2(_1172_),
    .B1(_1174_),
    .B2(\as2650.psu[3] ),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5020_ (.A1(_1188_),
    .A2(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5021_ (.A1(_1182_),
    .A2(_1134_),
    .B1(_3569_),
    .B2(_1183_),
    .C(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5022_ (.A1(\as2650.psu[0] ),
    .A2(_1175_),
    .B1(_0760_),
    .B2(\as2650.psu[5] ),
    .C(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5023_ (.A1(_0315_),
    .A2(_0261_),
    .A3(_1002_),
    .A4(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5024_ (.A1(_3134_),
    .A2(_0801_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5025_ (.A1(_1169_),
    .A2(_1181_),
    .B(_1193_),
    .C(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5026_ (.A1(_1160_),
    .A2(_0589_),
    .A3(_1194_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5027_ (.A1(_0803_),
    .A2(_1195_),
    .A3(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5028_ (.A1(_1161_),
    .A2(_1156_),
    .A3(_0804_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5029_ (.A1(_0584_),
    .A2(_1105_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5030_ (.A1(_0822_),
    .A2(_1198_),
    .B(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5031_ (.A1(_1053_),
    .A2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5032_ (.A1(_1121_),
    .A2(_0587_),
    .B(_1115_),
    .C(_1158_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5033_ (.A1(_1157_),
    .A2(_1159_),
    .B1(_1201_),
    .B2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5034_ (.I(_1093_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5035_ (.A1(_1152_),
    .A2(_1155_),
    .B1(_1203_),
    .B2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5036_ (.I0(_1205_),
    .I1(_1160_),
    .S(_1062_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5037_ (.A1(_1151_),
    .A2(_1206_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5038_ (.I(_1207_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5039_ (.I(_0888_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5040_ (.I(_0893_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5041_ (.I(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5042_ (.I(_0927_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5043_ (.I(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5044_ (.I(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5045_ (.A1(_0920_),
    .A2(_0926_),
    .B(_1213_),
    .C(_3264_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5046_ (.A1(_1210_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5047_ (.A1(_0899_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5048_ (.I(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5049_ (.I0(\as2650.stack[5][0] ),
    .I1(_1208_),
    .S(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5050_ (.I(_1218_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5051_ (.I(_0936_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5052_ (.I0(\as2650.stack[5][1] ),
    .I1(_1219_),
    .S(_1217_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_1220_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5054_ (.I0(\as2650.stack[5][2] ),
    .I1(_0942_),
    .S(_1217_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5055_ (.I(_1221_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5056_ (.I(_0947_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5057_ (.I0(\as2650.stack[5][3] ),
    .I1(_1222_),
    .S(_1217_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5058_ (.I(_1223_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5059_ (.I(\as2650.pc[4] ),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5060_ (.I(_1224_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5061_ (.I(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5062_ (.I(_1216_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5063_ (.I0(\as2650.stack[5][4] ),
    .I1(_1226_),
    .S(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5064_ (.I(_1228_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5065_ (.I(\as2650.pc[5] ),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5066_ (.I(_1229_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5067_ (.I0(\as2650.stack[5][5] ),
    .I1(_1230_),
    .S(_1227_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5068_ (.I(_1231_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5069_ (.I(_0964_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5070_ (.I0(\as2650.stack[5][6] ),
    .I1(_1232_),
    .S(_1227_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5071_ (.I(_1233_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5072_ (.I(_0969_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5074_ (.I0(\as2650.stack[5][7] ),
    .I1(_1235_),
    .S(_1227_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5075_ (.I(_1236_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5076_ (.I(_0976_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5077_ (.I(_1216_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5078_ (.I0(\as2650.stack[5][8] ),
    .I1(_1237_),
    .S(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5079_ (.I(_1239_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5080_ (.I(\as2650.pc[9] ),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5081_ (.I(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5082_ (.I0(\as2650.stack[5][9] ),
    .I1(_1241_),
    .S(_1238_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5083_ (.I(_1242_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5084_ (.I(\as2650.pc[10] ),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5085_ (.I(_1243_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5086_ (.I0(\as2650.stack[5][10] ),
    .I1(_1244_),
    .S(_1238_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5087_ (.I(_1245_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5088_ (.I(\as2650.pc[11] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5089_ (.I(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5090_ (.I0(\as2650.stack[5][11] ),
    .I1(_1247_),
    .S(_1238_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5091_ (.I(_1248_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5092_ (.I(\as2650.pc[12] ),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5093_ (.I0(\as2650.stack[5][12] ),
    .I1(_1249_),
    .S(_1216_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(_1250_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_0896_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5098_ (.A1(_1210_),
    .A2(_0930_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5099_ (.A1(_1253_),
    .A2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5100_ (.I(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5101_ (.I0(\as2650.stack[4][0] ),
    .I1(_1208_),
    .S(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5102_ (.I(_1257_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5103_ (.I0(\as2650.stack[4][1] ),
    .I1(_1219_),
    .S(_1256_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5104_ (.I(_1258_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5105_ (.I0(\as2650.stack[4][2] ),
    .I1(_0942_),
    .S(_1256_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5106_ (.I(_1259_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5107_ (.I0(\as2650.stack[4][3] ),
    .I1(_1222_),
    .S(_1256_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5108_ (.I(_1260_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5109_ (.I(_1255_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5110_ (.I0(\as2650.stack[4][4] ),
    .I1(_1226_),
    .S(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5111_ (.I(_1262_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5112_ (.I0(\as2650.stack[4][5] ),
    .I1(_1230_),
    .S(_1261_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5113_ (.I(_1263_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5114_ (.I0(\as2650.stack[4][6] ),
    .I1(_1232_),
    .S(_1261_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5115_ (.I(_1264_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5116_ (.I0(\as2650.stack[4][7] ),
    .I1(_1235_),
    .S(_1261_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5117_ (.I(_1265_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5118_ (.I(_1255_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5119_ (.I0(\as2650.stack[4][8] ),
    .I1(_1237_),
    .S(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5120_ (.I(_1267_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5121_ (.I0(\as2650.stack[4][9] ),
    .I1(_1241_),
    .S(_1266_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5122_ (.I(_1268_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5123_ (.I0(\as2650.stack[4][10] ),
    .I1(_1244_),
    .S(_1266_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5124_ (.I(_1269_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5125_ (.I0(\as2650.stack[4][11] ),
    .I1(_1247_),
    .S(_1266_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5126_ (.I(_1270_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5127_ (.I0(\as2650.stack[4][12] ),
    .I1(_1249_),
    .S(_1255_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5128_ (.I(_1271_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5129_ (.I(\as2650.stack_ptr[2] ),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5130_ (.A1(_1272_),
    .A2(_1253_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5131_ (.A1(_1214_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5132_ (.I(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5133_ (.I(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5134_ (.I(_1274_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5135_ (.A1(\as2650.stack[3][0] ),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5136_ (.A1(_0892_),
    .A2(_1276_),
    .B(_1278_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(\as2650.stack[3][1] ),
    .A2(_1277_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5138_ (.A1(_0939_),
    .A2(_1276_),
    .B(_1279_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(\as2650.stack[3][2] ),
    .A2(_1277_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5140_ (.A1(_0945_),
    .A2(_1276_),
    .B(_1280_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(\as2650.stack[3][3] ),
    .A2(_1277_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5142_ (.A1(_0951_),
    .A2(_1276_),
    .B(_1281_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5143_ (.I(_1275_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5144_ (.I(_1274_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5145_ (.A1(\as2650.stack[3][4] ),
    .A2(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5146_ (.A1(_0955_),
    .A2(_1282_),
    .B(_1284_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5147_ (.A1(\as2650.stack[3][5] ),
    .A2(_1283_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5148_ (.A1(_0962_),
    .A2(_1282_),
    .B(_1285_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(\as2650.stack[3][6] ),
    .A2(_1283_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5150_ (.A1(_0967_),
    .A2(_1282_),
    .B(_1286_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(\as2650.stack[3][7] ),
    .A2(_1283_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5152_ (.A1(_0972_),
    .A2(_1282_),
    .B(_1287_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5153_ (.I0(_0977_),
    .I1(\as2650.stack[3][8] ),
    .S(_1275_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5154_ (.I(_1288_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5155_ (.I(_1275_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5156_ (.I(_1274_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5157_ (.A1(\as2650.stack[3][9] ),
    .A2(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5158_ (.A1(_0981_),
    .A2(_1289_),
    .B(_1291_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(\as2650.stack[3][10] ),
    .A2(_1290_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5160_ (.A1(_0987_),
    .A2(_1289_),
    .B(_1292_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(\as2650.stack[3][11] ),
    .A2(_1290_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5162_ (.A1(_0991_),
    .A2(_1289_),
    .B(_1293_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(\as2650.stack[3][12] ),
    .A2(_1290_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5164_ (.A1(_0995_),
    .A2(_1289_),
    .B(_1294_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5165_ (.I(_3151_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5166_ (.I(_1032_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5167_ (.A1(_3180_),
    .A2(_0917_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5168_ (.A1(_0640_),
    .A2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5169_ (.I(_1298_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5170_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5171_ (.A1(_0588_),
    .A2(_0678_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5172_ (.A1(_0621_),
    .A2(_1300_),
    .B(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5173_ (.A1(_1295_),
    .A2(_3171_),
    .A3(_1296_),
    .A4(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5174_ (.I(_1303_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5175_ (.I(_1128_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5176_ (.A1(_0903_),
    .A2(_1033_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5177_ (.I(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5178_ (.A1(_1305_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5179_ (.I(_3199_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(_1296_),
    .A2(_1309_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5181_ (.A1(_1303_),
    .A2(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5182_ (.I(_1311_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5183_ (.A1(_1165_),
    .A2(_1304_),
    .B1(_1308_),
    .B2(_1312_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5184_ (.I(_1129_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5185_ (.A1(_1313_),
    .A2(_1307_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5186_ (.A1(_0826_),
    .A2(_1304_),
    .B1(_1312_),
    .B2(_1314_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5187_ (.A1(_0833_),
    .A2(_1304_),
    .B1(_1312_),
    .B2(_1130_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5188_ (.I(_1315_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5189_ (.A1(_0676_),
    .A2(_0922_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5190_ (.I(_1316_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5191_ (.I(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5192_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5193_ (.A1(_1319_),
    .A2(_1303_),
    .B(_0447_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5194_ (.I0(_1320_),
    .I1(_0873_),
    .S(_1311_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5195_ (.I(_1321_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5196_ (.I(_1109_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5197_ (.A1(_1025_),
    .A2(_1304_),
    .B1(_1312_),
    .B2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5198_ (.I(_1323_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5199_ (.I(_1137_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5200_ (.A1(_1026_),
    .A2(_1303_),
    .B1(_1311_),
    .B2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5201_ (.I(_1325_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(_0930_),
    .A2(_1273_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5203_ (.I(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5204_ (.I(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(_1326_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(\as2650.stack[2][0] ),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5207_ (.A1(_0892_),
    .A2(_1328_),
    .B(_1330_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5208_ (.A1(\as2650.stack[2][1] ),
    .A2(_1329_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5209_ (.A1(_0939_),
    .A2(_1328_),
    .B(_1331_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5210_ (.A1(\as2650.stack[2][2] ),
    .A2(_1329_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5211_ (.A1(_0945_),
    .A2(_1328_),
    .B(_1332_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5212_ (.A1(\as2650.stack[2][3] ),
    .A2(_1329_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5213_ (.A1(_0951_),
    .A2(_1328_),
    .B(_1333_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5214_ (.I(_1327_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5215_ (.I(_1326_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5216_ (.A1(\as2650.stack[2][4] ),
    .A2(_1335_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5217_ (.A1(_0955_),
    .A2(_1334_),
    .B(_1336_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5218_ (.A1(\as2650.stack[2][5] ),
    .A2(_1335_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5219_ (.A1(_0962_),
    .A2(_1334_),
    .B(_1337_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5220_ (.A1(\as2650.stack[2][6] ),
    .A2(_1335_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5221_ (.A1(_0967_),
    .A2(_1334_),
    .B(_1338_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(\as2650.stack[2][7] ),
    .A2(_1335_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5223_ (.A1(_0972_),
    .A2(_1334_),
    .B(_1339_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5224_ (.I0(_0977_),
    .I1(\as2650.stack[2][8] ),
    .S(_1327_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5225_ (.I(_1340_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5226_ (.I(_1327_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5227_ (.I(_1326_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5228_ (.A1(\as2650.stack[2][9] ),
    .A2(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5229_ (.A1(_0981_),
    .A2(_1341_),
    .B(_1343_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5230_ (.A1(\as2650.stack[2][10] ),
    .A2(_1342_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5231_ (.A1(_0987_),
    .A2(_1341_),
    .B(_1344_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(\as2650.stack[2][11] ),
    .A2(_1342_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5233_ (.A1(_0991_),
    .A2(_1341_),
    .B(_1345_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(\as2650.stack[2][12] ),
    .A2(_1342_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5235_ (.A1(_0995_),
    .A2(_1341_),
    .B(_1346_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5236_ (.A1(_0672_),
    .A2(_0682_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5237_ (.I(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5238_ (.I0(_0669_),
    .I1(\as2650.r123_2[1][0] ),
    .S(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5239_ (.I(_1349_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5240_ (.I(_1348_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5241_ (.I(_1348_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5242_ (.A1(\as2650.r123_2[1][1] ),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5243_ (.A1(_0706_),
    .A2(_1350_),
    .B(_1352_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_1351_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5245_ (.A1(_0723_),
    .A2(_1350_),
    .B(_1353_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5246_ (.I(_1347_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5247_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5248_ (.A1(_0737_),
    .A2(_1350_),
    .B(_1355_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_1354_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5250_ (.A1(_0754_),
    .A2(_1350_),
    .B(_1356_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5251_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_1354_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5252_ (.A1(_0770_),
    .A2(_1351_),
    .B(_1357_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5253_ (.I0(_0783_),
    .I1(\as2650.r123_2[1][6] ),
    .S(_1348_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5254_ (.I(_1358_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5255_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_1354_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5256_ (.A1(_0796_),
    .A2(_1351_),
    .B(_1359_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5257_ (.A1(_0895_),
    .A2(_1253_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_0930_),
    .A2(_1360_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5259_ (.I(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5260_ (.I(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5261_ (.I(_1361_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(\as2650.stack[0][0] ),
    .A2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5263_ (.A1(_0892_),
    .A2(_1363_),
    .B(_1365_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5264_ (.A1(\as2650.stack[0][1] ),
    .A2(_1364_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5265_ (.A1(_0939_),
    .A2(_1363_),
    .B(_1366_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(\as2650.stack[0][2] ),
    .A2(_1364_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5267_ (.A1(_0944_),
    .A2(_1363_),
    .B(_1367_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(\as2650.stack[0][3] ),
    .A2(_1364_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5269_ (.A1(_0950_),
    .A2(_1363_),
    .B(_1368_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5270_ (.I(_1362_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5271_ (.I(_1361_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5272_ (.A1(\as2650.stack[0][4] ),
    .A2(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5273_ (.A1(_0954_),
    .A2(_1369_),
    .B(_1371_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(\as2650.stack[0][5] ),
    .A2(_1370_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5275_ (.A1(_0961_),
    .A2(_1369_),
    .B(_1372_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5276_ (.A1(\as2650.stack[0][6] ),
    .A2(_1370_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5277_ (.A1(_0966_),
    .A2(_1369_),
    .B(_1373_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(\as2650.stack[0][7] ),
    .A2(_1370_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5279_ (.A1(_0971_),
    .A2(_1369_),
    .B(_1374_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5280_ (.I0(_0977_),
    .I1(\as2650.stack[0][8] ),
    .S(_1362_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5281_ (.I(_1375_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5282_ (.I(_1362_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5283_ (.I(_1361_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(\as2650.stack[0][9] ),
    .A2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5285_ (.A1(_0981_),
    .A2(_1376_),
    .B(_1378_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5286_ (.A1(\as2650.stack[0][10] ),
    .A2(_1377_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5287_ (.A1(_0986_),
    .A2(_1376_),
    .B(_1379_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5288_ (.A1(\as2650.stack[0][11] ),
    .A2(_1377_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5289_ (.A1(_0991_),
    .A2(_1376_),
    .B(_1380_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5290_ (.A1(\as2650.stack[0][12] ),
    .A2(_1377_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5291_ (.A1(_0995_),
    .A2(_1376_),
    .B(_1381_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5292_ (.A1(_1214_),
    .A2(_1360_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5293_ (.I(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5294_ (.I(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5295_ (.I(_1382_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(\as2650.stack[1][0] ),
    .A2(_1385_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5297_ (.A1(_0891_),
    .A2(_1384_),
    .B(_1386_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5298_ (.A1(\as2650.stack[1][1] ),
    .A2(_1385_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5299_ (.A1(_0938_),
    .A2(_1384_),
    .B(_1387_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5300_ (.A1(\as2650.stack[1][2] ),
    .A2(_1385_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5301_ (.A1(_0944_),
    .A2(_1384_),
    .B(_1388_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(\as2650.stack[1][3] ),
    .A2(_1385_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5303_ (.A1(_0950_),
    .A2(_1384_),
    .B(_1389_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5304_ (.I(_1383_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5305_ (.I(_1382_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5306_ (.A1(\as2650.stack[1][4] ),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5307_ (.A1(_0954_),
    .A2(_1390_),
    .B(_1392_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5308_ (.A1(\as2650.stack[1][5] ),
    .A2(_1391_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5309_ (.A1(_0961_),
    .A2(_1390_),
    .B(_1393_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(\as2650.stack[1][6] ),
    .A2(_1391_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5311_ (.A1(_0966_),
    .A2(_1390_),
    .B(_1394_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5312_ (.A1(\as2650.stack[1][7] ),
    .A2(_1391_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5313_ (.A1(_0971_),
    .A2(_1390_),
    .B(_1395_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5314_ (.I0(_1237_),
    .I1(\as2650.stack[1][8] ),
    .S(_1383_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5315_ (.I(_1396_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5316_ (.I(_1383_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5317_ (.I(_1382_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(\as2650.stack[1][9] ),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5319_ (.A1(_0980_),
    .A2(_1397_),
    .B(_1399_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5320_ (.A1(\as2650.stack[1][10] ),
    .A2(_1398_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5321_ (.A1(_0986_),
    .A2(_1397_),
    .B(_1400_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5322_ (.A1(\as2650.stack[1][11] ),
    .A2(_1398_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(_0990_),
    .A2(_1397_),
    .B(_1401_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5324_ (.A1(\as2650.stack[1][12] ),
    .A2(_1398_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5325_ (.A1(_0994_),
    .A2(_1397_),
    .B(_1402_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5326_ (.I(\as2650.r123[3][0] ),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5327_ (.I(_1403_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(\as2650.r123[3][1] ),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_1404_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5330_ (.I(\as2650.r123[3][2] ),
    .Z(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5331_ (.I(_1405_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5332_ (.I(\as2650.r123[3][3] ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5333_ (.I(_1406_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5334_ (.I(\as2650.r123[3][4] ),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5335_ (.I(_1407_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5336_ (.I(\as2650.r123[3][5] ),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5337_ (.I(_1408_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5338_ (.I(\as2650.r123[3][6] ),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5339_ (.I(_1409_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5340_ (.I(\as2650.r123[3][7] ),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5341_ (.I(_1410_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_0928_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_0675_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5344_ (.I(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5345_ (.I(_0903_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5346_ (.A1(_3197_),
    .A2(_0905_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(_1414_),
    .A2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5348_ (.A1(_0676_),
    .A2(_1297_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5349_ (.A1(_0817_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5350_ (.A1(_1107_),
    .A2(_1298_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5351_ (.I(_0316_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5352_ (.A1(_1420_),
    .A2(_0623_),
    .A3(_0917_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5353_ (.A1(_1416_),
    .A2(_1418_),
    .A3(_1419_),
    .B(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5354_ (.I(_3261_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5355_ (.I(_1006_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5356_ (.I(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5357_ (.I(_0925_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5358_ (.I(_1317_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5359_ (.I(_3209_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5360_ (.A1(_1428_),
    .A2(_0814_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5361_ (.A1(_1425_),
    .A2(_1426_),
    .B(_1427_),
    .C(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(_0677_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5363_ (.I(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_1051_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5365_ (.A1(_1412_),
    .A2(_1432_),
    .A3(_1433_),
    .A4(_0917_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5366_ (.A1(_1423_),
    .A2(_1430_),
    .A3(_1434_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5367_ (.I(_1424_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5368_ (.I(_0906_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5369_ (.I(_1417_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5370_ (.I(_3181_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5371_ (.I(_1439_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5372_ (.I(_0838_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5373_ (.I(_1317_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5374_ (.A1(_1440_),
    .A2(_1441_),
    .A3(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5375_ (.A1(_1436_),
    .A2(_1437_),
    .A3(_1438_),
    .A4(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5376_ (.A1(_3214_),
    .A2(_0919_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5377_ (.A1(_3349_),
    .A2(_0863_),
    .B1(_0915_),
    .B2(_1428_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5378_ (.I(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5379_ (.A1(_1444_),
    .A2(_1445_),
    .A3(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5380_ (.A1(_1413_),
    .A2(_1422_),
    .B(_1435_),
    .C(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5381_ (.I(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5382_ (.A1(_1411_),
    .A2(_1450_),
    .B(_0885_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5383_ (.A1(_1411_),
    .A2(_1450_),
    .B(_1451_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5384_ (.I(_1439_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5385_ (.I(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5386_ (.A1(\as2650.stack_ptr[1] ),
    .A2(\as2650.stack_ptr[0] ),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5387_ (.I(_1454_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5388_ (.A1(\as2650.stack_ptr[1] ),
    .A2(\as2650.stack_ptr[0] ),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5389_ (.A1(_1455_),
    .A2(_1456_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5390_ (.I(_1457_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5391_ (.A1(_1453_),
    .A2(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5392_ (.A1(_0899_),
    .A2(_1449_),
    .B(_0885_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5393_ (.A1(_1450_),
    .A2(_1459_),
    .B(_1460_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_0675_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5395_ (.I(_1461_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5396_ (.A1(_1462_),
    .A2(_1458_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5397_ (.A1(_1272_),
    .A2(_1454_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5398_ (.I(_1464_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5399_ (.A1(_0896_),
    .A2(_0927_),
    .B(\as2650.stack_ptr[2] ),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5400_ (.A1(_1465_),
    .A2(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5402_ (.I(_1468_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5403_ (.A1(_1463_),
    .A2(_1469_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5404_ (.A1(_0895_),
    .A2(_1449_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5405_ (.I(_3449_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5406_ (.I(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5407_ (.A1(_1450_),
    .A2(_1470_),
    .B(_1471_),
    .C(_1473_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5408_ (.A1(_0671_),
    .A2(_0682_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5409_ (.I(_1474_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5410_ (.I0(_0669_),
    .I1(\as2650.r123_2[0][0] ),
    .S(_1475_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_1476_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5412_ (.I(_1475_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5413_ (.I(_1475_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(\as2650.r123_2[0][1] ),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5415_ (.A1(_0706_),
    .A2(_1477_),
    .B(_1479_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(\as2650.r123_2[0][2] ),
    .A2(_1478_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5417_ (.A1(_0723_),
    .A2(_1477_),
    .B(_1480_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5418_ (.I(_1474_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5419_ (.A1(\as2650.r123_2[0][3] ),
    .A2(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5420_ (.A1(_0737_),
    .A2(_1477_),
    .B(_1482_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5421_ (.A1(\as2650.r123_2[0][4] ),
    .A2(_1481_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5422_ (.A1(_0754_),
    .A2(_1477_),
    .B(_1483_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5423_ (.A1(\as2650.r123_2[0][5] ),
    .A2(_1481_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5424_ (.A1(_0770_),
    .A2(_1478_),
    .B(_1484_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5425_ (.I0(_0783_),
    .I1(\as2650.r123_2[0][6] ),
    .S(_1475_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_1485_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_1481_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5428_ (.A1(_0796_),
    .A2(_1478_),
    .B(_1486_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5429_ (.I(_1175_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5430_ (.I(_3196_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5431_ (.A1(_3154_),
    .A2(_3279_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5432_ (.A1(_3195_),
    .A2(_1488_),
    .A3(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5433_ (.A1(_0906_),
    .A2(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5434_ (.I(_3239_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5435_ (.A1(\as2650.cycle[6] ),
    .A2(_3196_),
    .A3(_1489_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5436_ (.A1(_3305_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5437_ (.A1(_1492_),
    .A2(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5438_ (.A1(_1007_),
    .A2(_1491_),
    .A3(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5439_ (.A1(_0909_),
    .A2(_1496_),
    .B(_1082_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5440_ (.I(_0902_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5442_ (.I(_1316_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5443_ (.A1(_1045_),
    .A2(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5444_ (.I(_0655_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5445_ (.A1(_0810_),
    .A2(_1080_),
    .A3(_1000_),
    .A4(_0919_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5446_ (.A1(_3208_),
    .A2(_3194_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5447_ (.A1(_1504_),
    .A2(_0851_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5448_ (.A1(_0315_),
    .A2(_0318_),
    .B(_1299_),
    .C(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5449_ (.A1(_3264_),
    .A2(_1502_),
    .A3(_1503_),
    .A4(_1506_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5450_ (.I(_3278_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5451_ (.A1(_0835_),
    .A2(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5452_ (.A1(_1414_),
    .A2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5453_ (.I(_1510_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5454_ (.A1(_1439_),
    .A2(_0913_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5455_ (.A1(_0999_),
    .A2(_0924_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5456_ (.A1(_1511_),
    .A2(_1512_),
    .A3(_1416_),
    .A4(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5457_ (.I(\as2650.cycle[6] ),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5458_ (.A1(_1515_),
    .A2(_1490_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5459_ (.A1(_0999_),
    .A2(_1417_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5460_ (.A1(_3212_),
    .A2(_1416_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5461_ (.A1(_0901_),
    .A2(_1517_),
    .B(_1518_),
    .C(_1014_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5462_ (.A1(_1419_),
    .A2(_1514_),
    .B1(_1516_),
    .B2(_1081_),
    .C(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5463_ (.A1(_1499_),
    .A2(_1501_),
    .B(_1507_),
    .C(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5464_ (.A1(_1497_),
    .A2(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5465_ (.I(_1522_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5466_ (.I(_1523_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5467_ (.I(\as2650.addr_buff[0] ),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5468_ (.I(_1522_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5469_ (.A1(_1525_),
    .A2(_1526_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5470_ (.A1(_1487_),
    .A2(_1524_),
    .B(_1527_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(\as2650.addr_buff[1] ),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5472_ (.I(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5473_ (.I(_1522_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5474_ (.A1(_1529_),
    .A2(_1530_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5475_ (.A1(_1173_),
    .A2(_1524_),
    .B(_1531_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5476_ (.I(_3568_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5477_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5478_ (.I(_1533_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5479_ (.I(\as2650.addr_buff[2] ),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(_1535_),
    .A2(_1530_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5481_ (.A1(_1534_),
    .A2(_1524_),
    .B(_1536_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5482_ (.I(_1174_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5483_ (.I(\as2650.addr_buff[3] ),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5484_ (.A1(_1538_),
    .A2(_1530_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5485_ (.A1(_1537_),
    .A2(_1524_),
    .B(_1539_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5486_ (.I(_1184_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5487_ (.I(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5488_ (.I(\as2650.addr_buff[4] ),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(_1542_),
    .A2(_1530_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5490_ (.A1(_1541_),
    .A2(_1526_),
    .B(_1543_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5491_ (.I(_0760_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5492_ (.A1(_3233_),
    .A2(_1523_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5493_ (.A1(_1544_),
    .A2(_1526_),
    .B(_1545_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5494_ (.I(_1187_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5495_ (.A1(_3234_),
    .A2(_1523_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5496_ (.A1(_1546_),
    .A2(_1526_),
    .B(_1547_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5497_ (.I(_0316_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5498_ (.I0(_1324_),
    .I1(_1548_),
    .S(_1523_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_1549_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5500_ (.I(net24),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5501_ (.I(_1510_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5502_ (.A1(_3397_),
    .A2(_3221_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5503_ (.A1(_0837_),
    .A2(_1551_),
    .A3(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5504_ (.I(_1017_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5505_ (.A1(_1033_),
    .A2(_1045_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5506_ (.A1(_0646_),
    .A2(_0814_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5507_ (.A1(_3223_),
    .A2(_1556_),
    .B(_1504_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5508_ (.I(_0902_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5509_ (.A1(_0913_),
    .A2(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(_1557_),
    .A2(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5511_ (.A1(_1554_),
    .A2(_1555_),
    .A3(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5512_ (.I(_1108_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5513_ (.A1(_1562_),
    .A2(_1018_),
    .B(_1015_),
    .C(_3261_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5514_ (.A1(_1437_),
    .A2(_1008_),
    .B(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5515_ (.A1(_1553_),
    .A2(_1561_),
    .A3(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5516_ (.I(_1048_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5517_ (.I(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5518_ (.I(_1052_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5519_ (.A1(_1567_),
    .A2(_1568_),
    .B(_1518_),
    .C(_1565_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5520_ (.A1(_1550_),
    .A2(_1565_),
    .B(_1569_),
    .C(_1473_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5521_ (.I(_1036_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5522_ (.I(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5523_ (.I(_1428_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5524_ (.I(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5525_ (.A1(_1571_),
    .A2(_1573_),
    .A3(_0875_),
    .A4(_3221_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5526_ (.I(_0884_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5527_ (.A1(net22),
    .A2(_1574_),
    .B(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5528_ (.A1(_3479_),
    .A2(_1574_),
    .B(_1576_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5529_ (.A1(_3173_),
    .A2(_3279_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5530_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5531_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5532_ (.A1(_1452_),
    .A2(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5533_ (.A1(_0837_),
    .A2(_1043_),
    .B(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5534_ (.I(_1143_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5535_ (.A1(_1582_),
    .A2(_1035_),
    .B1(_0852_),
    .B2(_1556_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5536_ (.I(_1552_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5537_ (.A1(_3365_),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5538_ (.A1(_0850_),
    .A2(_1553_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5539_ (.A1(_1034_),
    .A2(_1013_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5540_ (.A1(_1036_),
    .A2(_1307_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5541_ (.A1(_1585_),
    .A2(_1586_),
    .A3(_1587_),
    .A4(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5542_ (.A1(_1581_),
    .A2(_1583_),
    .A3(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5543_ (.I(_1149_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5544_ (.A1(net23),
    .A2(_1590_),
    .B(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5545_ (.A1(_3175_),
    .A2(_1590_),
    .B(_1592_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5546_ (.A1(_3308_),
    .A2(_1496_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5547_ (.A1(_3260_),
    .A2(_1032_),
    .A3(_0902_),
    .A4(_1491_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5548_ (.A1(_3232_),
    .A2(_0409_),
    .A3(_1024_),
    .A4(_1029_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5549_ (.A1(_0851_),
    .A2(_1055_),
    .B1(_1555_),
    .B2(_3165_),
    .C(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5550_ (.A1(_1593_),
    .A2(_1594_),
    .B(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5551_ (.A1(_1301_),
    .A2(_1500_),
    .B(_1518_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5552_ (.A1(_0315_),
    .A2(_0817_),
    .B(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5553_ (.I(_1490_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5554_ (.A1(_1515_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5555_ (.A1(_1080_),
    .A2(_1578_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5556_ (.I(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5557_ (.A1(_1156_),
    .A2(_1601_),
    .A3(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5558_ (.A1(_1515_),
    .A2(_1488_),
    .A3(_1489_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5559_ (.A1(_3306_),
    .A2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5560_ (.A1(_1603_),
    .A2(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5561_ (.A1(_1310_),
    .A2(_1559_),
    .A3(_1604_),
    .A4(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5562_ (.I(_1502_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5563_ (.A1(_1048_),
    .A2(_1035_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5564_ (.A1(_1440_),
    .A2(_1609_),
    .A3(_1610_),
    .A4(_0918_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5565_ (.A1(_0317_),
    .A2(\as2650.addr_buff[7] ),
    .A3(_3307_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5566_ (.A1(_1494_),
    .A2(_1612_),
    .B(_3212_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5567_ (.A1(_1599_),
    .A2(_1608_),
    .A3(_1611_),
    .A4(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5568_ (.A1(_1597_),
    .A2(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5569_ (.A1(_0860_),
    .A2(_0916_),
    .B(_0861_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5570_ (.A1(_1445_),
    .A2(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5571_ (.A1(_1032_),
    .A2(_1045_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5572_ (.A1(_0806_),
    .A2(_0852_),
    .B1(_1500_),
    .B2(_1618_),
    .C(\as2650.halted ),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(_1502_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5574_ (.A1(_1620_),
    .A2(_1056_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5575_ (.A1(_1586_),
    .A2(_1617_),
    .A3(_1619_),
    .A4(_1621_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5576_ (.A1(_1585_),
    .A2(_1587_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5577_ (.A1(_0876_),
    .A2(_3319_),
    .B(_1037_),
    .C(_1623_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5578_ (.A1(_0874_),
    .A2(_0829_),
    .B(_1622_),
    .C(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5579_ (.A1(_3210_),
    .A2(_3188_),
    .A3(_3370_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5580_ (.A1(_3514_),
    .A2(_3567_),
    .A3(_0334_),
    .A4(_1626_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5581_ (.A1(_0381_),
    .A2(_0488_),
    .A3(_0591_),
    .A4(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(_0537_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5583_ (.I(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5584_ (.A1(_1445_),
    .A2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5585_ (.A1(_1615_),
    .A2(_1625_),
    .A3(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5586_ (.I(_0850_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5587_ (.I(_1633_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5588_ (.A1(_0875_),
    .A2(_1634_),
    .A3(_1018_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5589_ (.I(_3251_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5590_ (.A1(_1566_),
    .A2(_0907_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5591_ (.A1(net53),
    .A2(_1636_),
    .B(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_0924_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5593_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5594_ (.A1(_1043_),
    .A2(_1640_),
    .B(net53),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5595_ (.I(_1609_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5596_ (.I(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5597_ (.A1(_1638_),
    .A2(_1641_),
    .B(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(_1296_),
    .A2(_3279_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5599_ (.I(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5600_ (.I(_1646_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5601_ (.A1(_1635_),
    .A2(_1644_),
    .B(_1647_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5602_ (.A1(net53),
    .A2(_1632_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5603_ (.A1(_1632_),
    .A2(_1648_),
    .B(_1649_),
    .C(_1473_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5604_ (.I(_1149_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5605_ (.A1(_1445_),
    .A2(_1630_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_1097_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5607_ (.I(_1652_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5608_ (.A1(_1653_),
    .A2(_1555_),
    .B(_1595_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5609_ (.I(_1438_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5610_ (.A1(_1309_),
    .A2(_1005_),
    .B(_1568_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5611_ (.A1(_1298_),
    .A2(_1618_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5612_ (.A1(_3175_),
    .A2(_1508_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5613_ (.A1(_0923_),
    .A2(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5614_ (.A1(_1509_),
    .A2(_1657_),
    .A3(_1659_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5615_ (.A1(_1655_),
    .A2(_1656_),
    .B(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(_0810_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5617_ (.I(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5618_ (.I(_1297_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5619_ (.I(_1046_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5620_ (.A1(_1663_),
    .A2(_0819_),
    .A3(_1664_),
    .A4(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5621_ (.A1(_1654_),
    .A2(_1625_),
    .A3(_1661_),
    .A4(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5622_ (.A1(_1651_),
    .A2(_1667_),
    .B(net25),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5623_ (.A1(_1156_),
    .A2(_1318_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5624_ (.A1(_0910_),
    .A2(_0925_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(_1000_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5626_ (.A1(_1671_),
    .A2(_1442_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5627_ (.A1(net25),
    .A2(_0911_),
    .A3(_1670_),
    .A4(_1672_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5628_ (.A1(_1669_),
    .A2(_1673_),
    .B(_1440_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5629_ (.I(_0900_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(net25),
    .A2(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5631_ (.A1(_1412_),
    .A2(_1584_),
    .A3(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5632_ (.A1(_1143_),
    .A2(_1642_),
    .A3(_1674_),
    .A4(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5633_ (.A1(_0909_),
    .A2(_1676_),
    .B(_1083_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5634_ (.A1(_1310_),
    .A2(_1678_),
    .A3(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5635_ (.A1(_1647_),
    .A2(_1651_),
    .A3(_1667_),
    .A4(_1680_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5636_ (.A1(_1650_),
    .A2(_1668_),
    .A3(_1681_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_1492_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5638_ (.I(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5639_ (.A1(_1562_),
    .A2(_1610_),
    .A3(_1588_),
    .A4(_1607_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5640_ (.A1(_0913_),
    .A2(_0908_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5641_ (.A1(_3260_),
    .A2(_1516_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5642_ (.A1(_1014_),
    .A2(_1686_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5643_ (.A1(_3304_),
    .A2(_1416_),
    .B(_1685_),
    .C(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _5644_ (.A1(_1683_),
    .A2(_1594_),
    .B(_1684_),
    .C(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5645_ (.I(_1646_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5646_ (.A1(_3233_),
    .A2(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5647_ (.A1(_3299_),
    .A2(_1689_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5648_ (.A1(_1689_),
    .A2(_1691_),
    .B(_1692_),
    .C(_1473_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5649_ (.A1(_3234_),
    .A2(_1690_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5650_ (.A1(_3297_),
    .A2(_1689_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5651_ (.I(_1472_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5652_ (.A1(_1689_),
    .A2(_1693_),
    .B(_1694_),
    .C(_1695_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_0869_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5654_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(_3316_),
    .A2(_1609_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5656_ (.A1(_1487_),
    .A2(_1697_),
    .B(_1698_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5657_ (.I(_0409_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5658_ (.I(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5659_ (.A1(_1701_),
    .A2(_1636_),
    .A3(_1027_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5660_ (.A1(_1675_),
    .A2(_1029_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _5661_ (.A1(_0874_),
    .A2(_1702_),
    .B(_1703_),
    .C(_3265_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5662_ (.I(_1704_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5663_ (.I0(_1699_),
    .I1(_3407_),
    .S(_1705_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5664_ (.I(_1706_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_1105_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5666_ (.I(_1707_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5667_ (.A1(_3493_),
    .A2(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5668_ (.A1(_1173_),
    .A2(_1643_),
    .B(_1709_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5669_ (.I0(_1710_),
    .I1(_3460_),
    .S(_1705_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5670_ (.I(_1711_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(_1704_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5672_ (.I(_3554_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5673_ (.I(_0823_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5674_ (.A1(_1534_),
    .A2(_0822_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_1713_),
    .A2(_1714_),
    .B(_1715_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5676_ (.A1(_3580_),
    .A2(_1712_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5677_ (.A1(_1712_),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5678_ (.I(_1620_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5679_ (.I(_1718_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(_0725_),
    .A2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5681_ (.A1(_1537_),
    .A2(_1697_),
    .B(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5682_ (.I0(_1721_),
    .I1(_0287_),
    .S(_1705_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5683_ (.I(_1722_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5684_ (.A1(_0363_),
    .A2(_1719_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5685_ (.A1(_1541_),
    .A2(_1697_),
    .B(_1723_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5686_ (.I0(_1724_),
    .I1(_0396_),
    .S(_1705_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1725_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5688_ (.A1(_1544_),
    .A2(_1718_),
    .B(_0870_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5689_ (.I0(_1726_),
    .I1(_0440_),
    .S(_1704_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_1727_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5691_ (.I(_0536_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5692_ (.I(_0854_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5693_ (.A1(_1728_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5694_ (.A1(_1546_),
    .A2(_1714_),
    .B(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5695_ (.I0(_1731_),
    .I1(_0501_),
    .S(_1704_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5696_ (.I(_1732_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5697_ (.A1(_1324_),
    .A2(_1714_),
    .B(_1199_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5698_ (.A1(_0560_),
    .A2(_1712_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_1712_),
    .A2(_1733_),
    .B(_1734_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5700_ (.I(_1149_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5701_ (.I(_1735_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5702_ (.A1(_1736_),
    .A2(_1038_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5703_ (.I(_1570_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5704_ (.I(_1295_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5705_ (.I(_1511_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5707_ (.I(_1740_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5708_ (.I(_1601_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5709_ (.A1(_1137_),
    .A2(_1636_),
    .B(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5710_ (.A1(_0874_),
    .A2(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5711_ (.A1(_1738_),
    .A2(_3201_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5712_ (.A1(_3195_),
    .A2(_1488_),
    .A3(_3200_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5713_ (.I(_1746_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5714_ (.A1(_3202_),
    .A2(_3251_),
    .B(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5715_ (.A1(_1548_),
    .A2(_1636_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5716_ (.A1(_1748_),
    .A2(_1749_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5717_ (.I(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5718_ (.A1(_1741_),
    .A2(_1744_),
    .A3(_1745_),
    .A4(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5719_ (.I(_1461_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5720_ (.A1(_1753_),
    .A2(_1663_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5721_ (.I(_1093_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5722_ (.A1(_1696_),
    .A2(_1754_),
    .B(_0851_),
    .C(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5723_ (.I(_1588_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5724_ (.A1(_1738_),
    .A2(_1319_),
    .B1(_1752_),
    .B2(_1756_),
    .C(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5725_ (.I(_1566_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1499_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_1040_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5728_ (.A1(_1053_),
    .A2(_1056_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5729_ (.A1(_1761_),
    .A2(_0863_),
    .B1(_1762_),
    .B2(_1562_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5730_ (.A1(_1760_),
    .A2(_1584_),
    .B(_1763_),
    .C(_1738_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5731_ (.I(_1300_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5732_ (.A1(_3246_),
    .A2(_1616_),
    .A3(_1629_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5733_ (.I(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5734_ (.I(_0921_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5735_ (.A1(_1295_),
    .A2(_0839_),
    .A3(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5736_ (.A1(_1295_),
    .A2(_1508_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5737_ (.A1(_1426_),
    .A2(_1767_),
    .A3(_1769_),
    .B1(_1670_),
    .B2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5738_ (.A1(_1413_),
    .A2(_1765_),
    .A3(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5739_ (.A1(_1573_),
    .A2(_1764_),
    .B(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5740_ (.A1(_1759_),
    .A2(_1035_),
    .A3(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5741_ (.A1(_1737_),
    .A2(_1738_),
    .B1(_1758_),
    .B2(_1774_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5742_ (.A1(_1736_),
    .A2(_1775_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5743_ (.A1(_1737_),
    .A2(_0621_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5744_ (.A1(_3175_),
    .A2(_1309_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(_1765_),
    .A2(_1659_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_1427_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5747_ (.A1(_1761_),
    .A2(_1777_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5748_ (.A1(_1779_),
    .A2(_1766_),
    .B1(_1780_),
    .B2(_0907_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_1438_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5750_ (.A1(_1777_),
    .A2(_1778_),
    .B1(_1781_),
    .B2(_1782_),
    .C(_1453_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5751_ (.A1(_1642_),
    .A2(_0863_),
    .A3(_1762_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5752_ (.A1(_1453_),
    .A2(_1780_),
    .A3(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(_1094_),
    .A2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5754_ (.I(_1516_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5755_ (.I(_1787_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(_1751_),
    .A2(_1777_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5757_ (.A1(_1788_),
    .A2(_1789_),
    .B(_0907_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5758_ (.A1(_1708_),
    .A2(_1754_),
    .B1(_1744_),
    .B2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5759_ (.A1(_1783_),
    .A2(_1786_),
    .B1(_1791_),
    .B2(_1759_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(_1423_),
    .A2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5761_ (.I(_1735_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5762_ (.A1(_1776_),
    .A2(_1793_),
    .B(_1794_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5763_ (.I(_1737_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5764_ (.I(_1472_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5765_ (.A1(_3185_),
    .A2(_1577_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5766_ (.I(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5768_ (.I(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5769_ (.I(_1551_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5770_ (.A1(_0904_),
    .A2(_3227_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5771_ (.A1(_1801_),
    .A2(_1658_),
    .A3(_1802_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5772_ (.A1(_0910_),
    .A2(_1640_),
    .A3(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5773_ (.A1(_1801_),
    .A2(_1802_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5774_ (.A1(_1663_),
    .A2(_1568_),
    .B1(_1438_),
    .B2(_1805_),
    .C(_1318_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5775_ (.A1(_0819_),
    .A2(_1802_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5776_ (.A1(_1804_),
    .A2(_1806_),
    .B1(_1807_),
    .B2(_1319_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5777_ (.A1(_3228_),
    .A2(_0825_),
    .B(_1413_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5778_ (.I(_3229_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5779_ (.A1(_1810_),
    .A2(_1053_),
    .B(_1802_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_1424_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5781_ (.A1(_1675_),
    .A2(_1812_),
    .B(_1018_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5782_ (.A1(_1811_),
    .A2(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5783_ (.A1(_1573_),
    .A2(_1808_),
    .B1(_1809_),
    .B2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5784_ (.A1(_1022_),
    .A2(_3318_),
    .A3(_1144_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5785_ (.A1(_1029_),
    .A2(_1816_),
    .B(_1805_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5786_ (.I(_1603_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5787_ (.A1(_1800_),
    .A2(_1815_),
    .B1(_1817_),
    .B2(_1818_),
    .C(_1571_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5788_ (.A1(_1795_),
    .A2(_0904_),
    .B(_1796_),
    .C(_1819_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5789_ (.A1(_0447_),
    .A2(_1025_),
    .A3(_1026_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5790_ (.I(_1787_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5791_ (.A1(_3225_),
    .A2(_3226_),
    .A3(_3363_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5792_ (.A1(_0904_),
    .A2(_3227_),
    .B(_3277_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5793_ (.A1(_1822_),
    .A2(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5794_ (.A1(_1748_),
    .A2(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5795_ (.I(_1747_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5796_ (.I(_1826_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5797_ (.A1(_1548_),
    .A2(_1820_),
    .B(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5798_ (.A1(_1825_),
    .A2(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5799_ (.A1(_1324_),
    .A2(_1820_),
    .A3(_1821_),
    .B(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5800_ (.A1(_0909_),
    .A2(_0919_),
    .B(_1824_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5801_ (.A1(_1637_),
    .A2(_1830_),
    .B1(_1831_),
    .B2(_1567_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5802_ (.I(_1512_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5803_ (.A1(_1135_),
    .A2(_1000_),
    .A3(_1500_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5804_ (.A1(_1421_),
    .A2(_1834_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5805_ (.A1(_1833_),
    .A2(_1835_),
    .B(_1737_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5806_ (.A1(_1795_),
    .A2(_3277_),
    .B1(_1832_),
    .B2(_1836_),
    .C(_1796_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(\as2650.cycle[4] ),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5808_ (.A1(_1570_),
    .A2(_1822_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5809_ (.A1(_1837_),
    .A2(_1838_),
    .B(_1575_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5810_ (.A1(_1837_),
    .A2(_1838_),
    .B(_1839_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(_1837_),
    .A2(_1838_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5812_ (.A1(\as2650.cycle[5] ),
    .A2(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5813_ (.A1(_1736_),
    .A2(_1841_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5814_ (.I(_1515_),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(\as2650.cycle[5] ),
    .A2(_1837_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5816_ (.A1(_1822_),
    .A2(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(_1842_),
    .A2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5818_ (.A1(_1842_),
    .A2(_1844_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5819_ (.I(_1601_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5820_ (.A1(_3202_),
    .A2(_3241_),
    .A3(_1847_),
    .B(_1603_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5821_ (.A1(_1845_),
    .A2(_1846_),
    .A3(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5822_ (.I(_1572_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5823_ (.A1(_1850_),
    .A2(_0833_),
    .A3(_1719_),
    .A4(_1818_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5824_ (.A1(_1423_),
    .A2(_1604_),
    .A3(_1849_),
    .A4(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5825_ (.A1(_1423_),
    .A2(_1842_),
    .B(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5826_ (.A1(_1736_),
    .A2(_1853_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5827_ (.I(_1554_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5828_ (.I(_1747_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5829_ (.I(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5830_ (.I(_1742_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5831_ (.A1(_1708_),
    .A2(_1856_),
    .A3(_1857_),
    .B(_1818_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5832_ (.A1(_3306_),
    .A2(_1845_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5833_ (.A1(_1854_),
    .A2(_1580_),
    .B1(_1858_),
    .B2(_1859_),
    .C(_1571_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5834_ (.A1(_1795_),
    .A2(_3306_),
    .B(_1796_),
    .C(_1860_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5835_ (.A1(_0853_),
    .A2(_0831_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5836_ (.A1(_1719_),
    .A2(_1003_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5837_ (.A1(_1861_),
    .A2(_1862_),
    .B(net4),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5838_ (.A1(\as2650.psu[7] ),
    .A2(_1157_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5839_ (.A1(_0826_),
    .A2(_1157_),
    .B(_1708_),
    .C(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5840_ (.A1(_0831_),
    .A2(_1199_),
    .B1(_1865_),
    .B2(_1003_),
    .C(_1571_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5841_ (.A1(_1182_),
    .A2(_1795_),
    .B1(_1863_),
    .B2(_1866_),
    .C(_1796_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5842_ (.A1(_1309_),
    .A2(_1508_),
    .B1(_1558_),
    .B2(_1420_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5843_ (.A1(_1107_),
    .A2(_0813_),
    .A3(_0852_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_0922_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5845_ (.A1(_1511_),
    .A2(_1437_),
    .A3(_1869_),
    .A4(_1618_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5846_ (.A1(_1417_),
    .A2(_1867_),
    .B(_1868_),
    .C(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5847_ (.A1(_0675_),
    .A2(_0821_),
    .A3(_0862_),
    .B(_1834_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5848_ (.I(_1594_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5849_ (.A1(_0843_),
    .A2(_0846_),
    .B(_3246_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5850_ (.A1(_1873_),
    .A2(_1660_),
    .A3(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5851_ (.A1(_1688_),
    .A2(_1871_),
    .A3(_1872_),
    .A4(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5852_ (.A1(_1165_),
    .A2(_0845_),
    .B(_0828_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5853_ (.A1(_3214_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5854_ (.A1(_1042_),
    .A2(_1033_),
    .B1(_1019_),
    .B2(_1797_),
    .C(_1306_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5855_ (.A1(_1878_),
    .A2(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5856_ (.A1(_3246_),
    .A2(_1024_),
    .B(_1037_),
    .C(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5857_ (.A1(_1619_),
    .A2(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5858_ (.A1(_1833_),
    .A2(_1422_),
    .B(_1596_),
    .C(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5859_ (.A1(_1876_),
    .A2(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5860_ (.I(_1884_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5861_ (.I(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5862_ (.A1(_1048_),
    .A2(_1645_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5863_ (.I(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5864_ (.I(_1885_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5865_ (.A1(_0890_),
    .A2(_1888_),
    .B(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5866_ (.A1(_0889_),
    .A2(_1432_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5867_ (.A1(_1616_),
    .A2(_1630_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5868_ (.A1(_3247_),
    .A2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5869_ (.I(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5870_ (.A1(_1441_),
    .A2(_0925_),
    .B(_1767_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5871_ (.I(_1895_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5872_ (.A1(_1640_),
    .A2(_1891_),
    .A3(_1894_),
    .B1(_1896_),
    .B2(_0890_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5873_ (.A1(_0888_),
    .A2(_3373_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5874_ (.A1(_1108_),
    .A2(_1442_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5875_ (.I(_1899_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5876_ (.A1(_1502_),
    .A2(_1317_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5877_ (.I(_1901_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5878_ (.I(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5879_ (.A1(_1898_),
    .A2(_1900_),
    .B1(_1903_),
    .B2(_0889_),
    .C(_1462_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5880_ (.A1(_0888_),
    .A2(_1432_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5881_ (.A1(_0833_),
    .A2(_1898_),
    .B(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5882_ (.I(_3373_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5883_ (.I(_1510_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5884_ (.A1(_1907_),
    .A2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5885_ (.A1(_1433_),
    .A2(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5886_ (.A1(_1525_),
    .A2(_0750_),
    .B(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5887_ (.A1(_0819_),
    .A2(_1906_),
    .B(_1911_),
    .C(_1655_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5888_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_3328_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5889_ (.A1(_1487_),
    .A2(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5890_ (.A1(_1907_),
    .A2(_1908_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5891_ (.A1(_1436_),
    .A2(_1914_),
    .B(_1915_),
    .C(_1517_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5892_ (.A1(_1912_),
    .A2(_1916_),
    .B(_1419_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5893_ (.A1(_1765_),
    .A2(_1897_),
    .B(_1904_),
    .C(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5894_ (.I(_1456_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_1919_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5896_ (.I(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5897_ (.I(_1466_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5898_ (.A1(\as2650.stack[7][0] ),
    .A2(_1465_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5899_ (.A1(_0898_),
    .A2(\as2650.stack[5][0] ),
    .B1(\as2650.stack[4][0] ),
    .B2(_0929_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5900_ (.A1(_1921_),
    .A2(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5901_ (.A1(\as2650.stack[6][0] ),
    .A2(_1921_),
    .B1(_1922_),
    .B2(_1923_),
    .C(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1013_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5903_ (.A1(_1253_),
    .A2(\as2650.stack[1][0] ),
    .B1(\as2650.stack[0][0] ),
    .B2(_1411_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5904_ (.I(_1919_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5905_ (.I(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5906_ (.A1(_0894_),
    .A2(\as2650.stack[3][0] ),
    .B1(\as2650.stack[2][0] ),
    .B2(_1930_),
    .C(_1469_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5907_ (.A1(_1921_),
    .A2(_1928_),
    .B(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5908_ (.A1(_1927_),
    .A2(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5909_ (.A1(_1208_),
    .A2(_1010_),
    .B1(_1926_),
    .B2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5910_ (.A1(_1918_),
    .A2(_1934_),
    .B(_1800_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5911_ (.A1(_0891_),
    .A2(_1886_),
    .B1(_1890_),
    .B2(_1935_),
    .C(_1591_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5912_ (.I(_1889_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5913_ (.A1(_0936_),
    .A2(_0887_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5914_ (.I(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5915_ (.I(_1887_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5916_ (.I(_1442_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5917_ (.A1(_0887_),
    .A2(\as2650.ins_reg[2] ),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5918_ (.A1(_0936_),
    .A2(_1941_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5919_ (.A1(_0868_),
    .A2(_1937_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5920_ (.A1(_1892_),
    .A2(_1942_),
    .B1(_1943_),
    .B2(_1893_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5921_ (.I(_1558_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5922_ (.A1(_1498_),
    .A2(_1051_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5923_ (.A1(_3507_),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_1528_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5924_ (.I(_0810_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5925_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5926_ (.A1(\as2650.pc[1] ),
    .A2(net6),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5927_ (.A1(_1949_),
    .A2(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5928_ (.A1(_1662_),
    .A2(_1951_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5929_ (.A1(_1948_),
    .A2(_1938_),
    .B(_1952_),
    .C(_1051_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5930_ (.A1(_1947_),
    .A2(_1953_),
    .B(_1620_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5931_ (.A1(_3371_),
    .A2(_1913_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5932_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_3138_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5933_ (.A1(_1171_),
    .A2(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5934_ (.A1(_1955_),
    .A2(_1957_),
    .B(_1558_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5935_ (.A1(_1955_),
    .A2(_1957_),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5936_ (.A1(_3506_),
    .A2(_1511_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5937_ (.A1(_0900_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5938_ (.A1(_1040_),
    .A2(_1938_),
    .B1(_1959_),
    .B2(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5939_ (.A1(_1639_),
    .A2(_1943_),
    .A3(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5940_ (.A1(_1639_),
    .A2(_1944_),
    .A3(_1954_),
    .B(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5941_ (.A1(_1609_),
    .A2(_1951_),
    .B(_1943_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5942_ (.A1(_1318_),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5943_ (.A1(_1940_),
    .A2(_1964_),
    .B(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5944_ (.A1(_1464_),
    .A2(_1466_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5945_ (.I(_1968_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5946_ (.I0(\as2650.stack[7][1] ),
    .I1(\as2650.stack[4][1] ),
    .I2(\as2650.stack[5][1] ),
    .I3(\as2650.stack[6][1] ),
    .S0(_0928_),
    .S1(_0897_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(_1919_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5948_ (.I(_0927_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5949_ (.A1(_0897_),
    .A2(\as2650.stack[1][1] ),
    .B1(\as2650.stack[0][1] ),
    .B2(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_1456_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5951_ (.A1(_0893_),
    .A2(\as2650.stack[3][1] ),
    .B1(\as2650.stack[2][1] ),
    .B2(_1974_),
    .C(_1467_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5952_ (.A1(_1971_),
    .A2(_1973_),
    .B(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5953_ (.A1(_1969_),
    .A2(_1970_),
    .B(_1976_),
    .C(_1927_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5954_ (.I(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5955_ (.A1(_1429_),
    .A2(_1938_),
    .B1(_1967_),
    .B2(_1462_),
    .C(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5956_ (.A1(_1939_),
    .A2(_1979_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5957_ (.I(_1884_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5958_ (.A1(_1888_),
    .A2(_1938_),
    .B(_1980_),
    .C(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5959_ (.A1(_0938_),
    .A2(_1936_),
    .B(_1982_),
    .C(_1695_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_1889_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5961_ (.I(_1885_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5962_ (.A1(_0941_),
    .A2(\as2650.pc[1] ),
    .A3(_0887_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5963_ (.A1(_0937_),
    .A2(_0889_),
    .B(_0943_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5964_ (.A1(_1985_),
    .A2(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5965_ (.I(_1896_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5966_ (.I(_1901_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5967_ (.A1(\as2650.pc[2] ),
    .A2(net7),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5968_ (.A1(\as2650.pc[1] ),
    .A2(_3505_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5969_ (.A1(_1949_),
    .A2(_1950_),
    .B(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5970_ (.A1(_1990_),
    .A2(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5971_ (.I(_1899_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5972_ (.A1(_1989_),
    .A2(_1987_),
    .B1(_1993_),
    .B2(_1994_),
    .C(_1753_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5973_ (.I(_1798_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5974_ (.A1(_1988_),
    .A2(_1995_),
    .B(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5975_ (.A1(_0711_),
    .A2(_1739_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5976_ (.A1(_3505_),
    .A2(_1956_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5977_ (.A1(_1955_),
    .A2(_1957_),
    .B(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5978_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_3328_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5979_ (.A1(_3568_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5980_ (.A1(_2000_),
    .A2(_2002_),
    .B(_0750_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5981_ (.A1(_2000_),
    .A2(_2002_),
    .B(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(_3156_),
    .A2(_0924_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5983_ (.I(_2005_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5984_ (.A1(_2004_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5985_ (.I(_1427_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5986_ (.A1(_1616_),
    .A2(_1630_),
    .B(_1108_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5987_ (.A1(_0937_),
    .A2(_1941_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5988_ (.A1(_0943_),
    .A2(_2010_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5989_ (.A1(_1431_),
    .A2(_1993_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5990_ (.A1(_1948_),
    .A2(_1987_),
    .B(_1671_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5991_ (.A1(\as2650.addr_buff[2] ),
    .A2(_1551_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5992_ (.A1(_0711_),
    .A2(_0921_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5993_ (.A1(_0818_),
    .A2(_2014_),
    .A3(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5994_ (.A1(_2012_),
    .A2(_2013_),
    .B(_2016_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5995_ (.I(_0821_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5996_ (.A1(_2009_),
    .A2(_2011_),
    .B1(_2017_),
    .B2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5997_ (.A1(_1297_),
    .A2(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5998_ (.A1(_1998_),
    .A2(_2007_),
    .B(_2008_),
    .C(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5999_ (.A1(\as2650.stack[7][2] ),
    .A2(_1465_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_1974_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6001_ (.I(_1251_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6002_ (.I(_1211_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6003_ (.A1(_2024_),
    .A2(\as2650.stack[5][2] ),
    .B1(\as2650.stack[4][2] ),
    .B2(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6004_ (.A1(_2023_),
    .A2(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6005_ (.A1(\as2650.stack[6][2] ),
    .A2(_1930_),
    .B1(_1922_),
    .B2(_2022_),
    .C(_2027_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6006_ (.A1(_2024_),
    .A2(\as2650.stack[1][2] ),
    .B1(\as2650.stack[0][2] ),
    .B2(_2025_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6007_ (.A1(_2023_),
    .A2(_2029_),
    .B(_1969_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6008_ (.A1(_1210_),
    .A2(\as2650.stack[3][2] ),
    .B1(\as2650.stack[2][2] ),
    .B2(_1930_),
    .C(_2030_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6009_ (.A1(_0867_),
    .A2(_2028_),
    .A3(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6010_ (.I(_0824_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6011_ (.I(_1440_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6012_ (.A1(_2033_),
    .A2(_1987_),
    .B(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6013_ (.A1(_1995_),
    .A2(_2021_),
    .B1(_2032_),
    .B2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1799_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6015_ (.A1(_1987_),
    .A2(_1997_),
    .B1(_2036_),
    .B2(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6016_ (.A1(_1984_),
    .A2(_2038_),
    .B(_1575_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6017_ (.A1(_0945_),
    .A2(_1983_),
    .B(_2039_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6018_ (.A1(_0947_),
    .A2(_1985_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6019_ (.A1(_3247_),
    .A2(_1299_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6020_ (.A1(_0947_),
    .A2(_0337_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6021_ (.A1(_0941_),
    .A2(net7),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6022_ (.I(_2043_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6023_ (.A1(_1990_),
    .A2(_1992_),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6024_ (.A1(_2042_),
    .A2(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6025_ (.A1(_2041_),
    .A2(_2046_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6026_ (.I(_1461_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6027_ (.A1(_1989_),
    .A2(_2040_),
    .B(_2047_),
    .C(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6028_ (.A1(_1988_),
    .A2(_2049_),
    .B(_1996_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6029_ (.A1(_0941_),
    .A2(_2010_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6030_ (.A1(_0949_),
    .A2(_2051_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6031_ (.I(_0857_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6032_ (.A1(_0832_),
    .A2(_2040_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6033_ (.A1(_2053_),
    .A2(_2046_),
    .B(_2054_),
    .C(_1433_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6034_ (.A1(_1132_),
    .A2(_1499_),
    .B1(_1946_),
    .B2(_1538_),
    .C(_1620_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6035_ (.A1(_2055_),
    .A2(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6036_ (.A1(_1894_),
    .A2(_2052_),
    .B(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6037_ (.I(_1908_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6038_ (.I(_2005_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6039_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_3140_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6040_ (.A1(_3568_),
    .A2(_2001_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6041_ (.A1(_2000_),
    .A2(_2002_),
    .B(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6042_ (.A1(_0338_),
    .A2(_2061_),
    .A3(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6043_ (.A1(_1425_),
    .A2(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6044_ (.A1(_1132_),
    .A2(_2059_),
    .B(_2060_),
    .C(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6045_ (.A1(_1869_),
    .A2(_2058_),
    .B(_2066_),
    .C(_2008_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6046_ (.A1(_2024_),
    .A2(\as2650.stack[5][3] ),
    .B1(\as2650.stack[4][3] ),
    .B2(_2025_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(\as2650.stack[7][3] ),
    .A2(_1922_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6048_ (.A1(_2023_),
    .A2(_2068_),
    .B(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6049_ (.A1(\as2650.stack[6][3] ),
    .A2(_1921_),
    .B(_1969_),
    .C(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6050_ (.I(_0896_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6051_ (.A1(_2072_),
    .A2(\as2650.stack[1][3] ),
    .B1(\as2650.stack[0][3] ),
    .B2(_1212_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6052_ (.I(_1968_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6053_ (.A1(_2023_),
    .A2(_2073_),
    .B(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6054_ (.A1(_1210_),
    .A2(\as2650.stack[3][3] ),
    .B1(\as2650.stack[2][3] ),
    .B2(_1930_),
    .C(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6055_ (.A1(_0866_),
    .A2(_2071_),
    .A3(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6056_ (.A1(_2033_),
    .A2(_2040_),
    .B(_2034_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6057_ (.A1(_2049_),
    .A2(_2067_),
    .B1(_2077_),
    .B2(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6058_ (.A1(_2040_),
    .A2(_2050_),
    .B1(_2079_),
    .B2(_2037_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6059_ (.A1(_1984_),
    .A2(_2080_),
    .B(_1575_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6060_ (.A1(_0951_),
    .A2(_1983_),
    .B(_2081_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6061_ (.A1(_0949_),
    .A2(_1985_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6062_ (.A1(_1225_),
    .A2(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6063_ (.I(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6064_ (.A1(_0953_),
    .A2(net9),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6065_ (.I(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(\as2650.pc[3] ),
    .A2(_0335_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6067_ (.A1(\as2650.pc[3] ),
    .A2(net8),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6068_ (.A1(_2088_),
    .A2(_2045_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6069_ (.A1(_2087_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6070_ (.A1(_2086_),
    .A2(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6071_ (.A1(_1902_),
    .A2(_2084_),
    .B1(_2091_),
    .B2(_1994_),
    .C(_1753_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6072_ (.A1(_1988_),
    .A2(_2092_),
    .B(_1996_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6073_ (.A1(_0948_),
    .A2(_2051_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6074_ (.A1(_1225_),
    .A2(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6075_ (.A1(_1125_),
    .A2(_1812_),
    .B1(_1007_),
    .B2(_1542_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6076_ (.A1(_1431_),
    .A2(_2091_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6077_ (.A1(_2053_),
    .A2(_2083_),
    .B(_2097_),
    .C(_1810_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6078_ (.A1(_2096_),
    .A2(_2098_),
    .B(_2018_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6079_ (.A1(_1894_),
    .A2(_2095_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6080_ (.A1(_0335_),
    .A2(_2061_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6081_ (.A1(_0335_),
    .A2(_2061_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6082_ (.A1(_2063_),
    .A2(_2101_),
    .B(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6083_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_3140_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6084_ (.A1(net9),
    .A2(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6085_ (.A1(_2103_),
    .A2(_2105_),
    .B(_0624_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6086_ (.A1(_2103_),
    .A2(_2105_),
    .B(_2106_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6087_ (.A1(_1125_),
    .A2(_2059_),
    .B(_2005_),
    .C(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6088_ (.A1(_1782_),
    .A2(_2100_),
    .B(_2108_),
    .C(_2008_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6089_ (.I(_1974_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6090_ (.I(_1251_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(_1211_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6092_ (.A1(_2111_),
    .A2(\as2650.stack[5][4] ),
    .B1(\as2650.stack[4][4] ),
    .B2(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6093_ (.A1(_2110_),
    .A2(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6094_ (.I(_1455_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6095_ (.A1(\as2650.stack[7][4] ),
    .A2(_2115_),
    .B1(_1971_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6096_ (.A1(_1469_),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6097_ (.A1(_2024_),
    .A2(\as2650.stack[1][4] ),
    .B1(\as2650.stack[0][4] ),
    .B2(_2025_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6098_ (.I(_0893_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6099_ (.A1(_2119_),
    .A2(\as2650.stack[3][4] ),
    .B1(\as2650.stack[2][4] ),
    .B2(_1929_),
    .C(_1468_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6100_ (.A1(_2110_),
    .A2(_2118_),
    .B(_2120_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_0814_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6102_ (.A1(_2114_),
    .A2(_2117_),
    .B(_2121_),
    .C(_2122_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6103_ (.A1(_2033_),
    .A2(_2084_),
    .B(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6104_ (.A1(_2092_),
    .A2(_2109_),
    .B1(_2124_),
    .B2(_1850_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6105_ (.A1(_2084_),
    .A2(_2093_),
    .B1(_2125_),
    .B2(_2037_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6106_ (.I(_0883_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6107_ (.A1(_1984_),
    .A2(_2126_),
    .B(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6108_ (.A1(_0955_),
    .A2(_1983_),
    .B(_2128_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_1885_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6110_ (.A1(_0953_),
    .A2(_0948_),
    .A3(_1985_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6111_ (.A1(_0960_),
    .A2(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6112_ (.A1(_0959_),
    .A2(net1),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6113_ (.I(_2132_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6114_ (.A1(_1224_),
    .A2(_0377_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6115_ (.A1(_2085_),
    .A2(_2090_),
    .B(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6116_ (.A1(_2133_),
    .A2(_2135_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6117_ (.A1(_1903_),
    .A2(_2131_),
    .B1(_2136_),
    .B2(_1900_),
    .C(_2048_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6118_ (.A1(_1988_),
    .A2(_2137_),
    .B(_1996_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6119_ (.I(_1945_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6120_ (.A1(_0375_),
    .A2(_2104_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6121_ (.A1(_2103_),
    .A2(_2105_),
    .B(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6122_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_3140_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6123_ (.A1(_0759_),
    .A2(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6124_ (.A1(_2141_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6125_ (.A1(_2141_),
    .A2(_2143_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6126_ (.A1(_2139_),
    .A2(_2144_),
    .A3(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6127_ (.A1(_0872_),
    .A2(_1740_),
    .B(_2006_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6128_ (.A1(_1229_),
    .A2(_1224_),
    .A3(_2094_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6129_ (.A1(_1225_),
    .A2(_2094_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6130_ (.A1(_0960_),
    .A2(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_2148_),
    .A2(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_1948_),
    .A2(_2136_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6133_ (.A1(_0832_),
    .A2(_2131_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6134_ (.A1(_1433_),
    .A2(_2152_),
    .A3(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6135_ (.A1(_0871_),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_3233_),
    .C(_1105_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6136_ (.A1(_2009_),
    .A2(_2151_),
    .B1(_2154_),
    .B2(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6137_ (.A1(_1664_),
    .A2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6138_ (.A1(_2146_),
    .A2(_2147_),
    .B(_1779_),
    .C(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6139_ (.I(_2074_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6140_ (.I0(\as2650.stack[7][5] ),
    .I1(\as2650.stack[4][5] ),
    .I2(\as2650.stack[5][5] ),
    .I3(\as2650.stack[6][5] ),
    .S0(_1972_),
    .S1(_2111_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6141_ (.A1(_2111_),
    .A2(\as2650.stack[1][5] ),
    .B1(\as2650.stack[0][5] ),
    .B2(_0929_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6142_ (.I(_1467_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6143_ (.A1(_1209_),
    .A2(\as2650.stack[3][5] ),
    .B1(\as2650.stack[2][5] ),
    .B2(_1920_),
    .C(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6144_ (.A1(_2110_),
    .A2(_2161_),
    .B(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6145_ (.A1(_2159_),
    .A2(_2160_),
    .B(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6146_ (.A1(_1429_),
    .A2(_2131_),
    .B1(_2165_),
    .B2(_1927_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6147_ (.A1(_2137_),
    .A2(_2158_),
    .B(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6148_ (.A1(_2131_),
    .A2(_2138_),
    .B1(_2167_),
    .B2(_2037_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6149_ (.A1(_2129_),
    .A2(_2168_),
    .B(_2127_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6150_ (.A1(_0962_),
    .A2(_1983_),
    .B(_2169_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6151_ (.A1(_1229_),
    .A2(_2130_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6152_ (.A1(_0964_),
    .A2(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6153_ (.I(_1896_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6154_ (.A1(\as2650.pc[6] ),
    .A2(net2),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6155_ (.A1(_1224_),
    .A2(net9),
    .B1(net1),
    .B2(\as2650.pc[5] ),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6156_ (.A1(_0960_),
    .A2(_0759_),
    .B(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6157_ (.I(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6158_ (.A1(_2085_),
    .A2(_2090_),
    .A3(_2133_),
    .B(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6159_ (.A1(_2173_),
    .A2(_2177_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6160_ (.A1(_1989_),
    .A2(_2171_),
    .B1(_2178_),
    .B2(_1994_),
    .C(_2048_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(_1798_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6162_ (.A1(_2172_),
    .A2(_2179_),
    .B(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6163_ (.A1(_0965_),
    .A2(_2148_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6164_ (.A1(_1662_),
    .A2(_2178_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_1431_),
    .A2(_2171_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6166_ (.A1(_1052_),
    .A2(_2183_),
    .A3(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6167_ (.A1(_1187_),
    .A2(_1812_),
    .B1(_1007_),
    .B2(_3387_),
    .C(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6168_ (.A1(_1894_),
    .A2(_2182_),
    .B1(_2186_),
    .B2(_1718_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6169_ (.A1(_0489_),
    .A2(_2142_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6170_ (.A1(_2141_),
    .A2(_2143_),
    .B(_2188_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6171_ (.A1(_0538_),
    .A2(_0473_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6172_ (.A1(_2189_),
    .A2(_2190_),
    .B(_0750_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6173_ (.A1(_2189_),
    .A2(_2190_),
    .B(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6174_ (.A1(_1322_),
    .A2(_2059_),
    .B(_2060_),
    .C(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6175_ (.A1(_1782_),
    .A2(_2187_),
    .B(_2193_),
    .C(_1779_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_1929_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6177_ (.A1(_2072_),
    .A2(\as2650.stack[1][6] ),
    .B1(\as2650.stack[0][6] ),
    .B2(_1972_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6178_ (.A1(_1971_),
    .A2(_2196_),
    .B(_2074_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6179_ (.A1(_0894_),
    .A2(\as2650.stack[3][6] ),
    .B1(\as2650.stack[2][6] ),
    .B2(_2195_),
    .C(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6180_ (.I(_1211_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6181_ (.A1(_2111_),
    .A2(\as2650.stack[5][6] ),
    .B1(\as2650.stack[4][6] ),
    .B2(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6182_ (.A1(\as2650.stack[7][6] ),
    .A2(_2115_),
    .B1(_1971_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6183_ (.A1(_2110_),
    .A2(_2200_),
    .B(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6184_ (.A1(_2159_),
    .A2(_2202_),
    .B(_2122_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6185_ (.A1(_2033_),
    .A2(_2171_),
    .B1(_2198_),
    .B2(_2203_),
    .C(_1452_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6186_ (.A1(_2179_),
    .A2(_2194_),
    .B(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6187_ (.I(_1799_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6188_ (.A1(_2171_),
    .A2(_2181_),
    .B1(_2205_),
    .B2(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6189_ (.A1(_2129_),
    .A2(_2207_),
    .B(_2127_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6190_ (.A1(_0967_),
    .A2(_1936_),
    .B(_2208_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6191_ (.A1(\as2650.pc[6] ),
    .A2(_1229_),
    .A3(_2130_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6192_ (.A1(_1234_),
    .A2(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6193_ (.I(_2041_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6194_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6195_ (.A1(\as2650.pc[6] ),
    .A2(_1185_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6196_ (.A1(_2173_),
    .A2(_2177_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6197_ (.A1(_2213_),
    .A2(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6198_ (.A1(_2212_),
    .A2(_2215_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6199_ (.A1(_2211_),
    .A2(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6200_ (.A1(_1903_),
    .A2(_2210_),
    .B(_2048_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6201_ (.A1(_1896_),
    .A2(_2217_),
    .A3(_2218_),
    .B(_2180_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_1893_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6203_ (.A1(_0965_),
    .A2(_2148_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6204_ (.A1(_1234_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(_1548_),
    .A2(_1908_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6206_ (.A1(_1136_),
    .A2(_0921_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6207_ (.A1(_0818_),
    .A2(_2223_),
    .A3(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6208_ (.A1(_1662_),
    .A2(_2216_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6209_ (.A1(_1948_),
    .A2(_2210_),
    .B(_2226_),
    .C(_1671_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6210_ (.A1(_2225_),
    .A2(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6211_ (.A1(_2220_),
    .A2(_2222_),
    .B1(_2228_),
    .B2(_1707_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6212_ (.I(_1185_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6213_ (.A1(_2230_),
    .A2(_0473_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6214_ (.A1(_2189_),
    .A2(_2190_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6215_ (.A1(_1135_),
    .A2(_3341_),
    .A3(_2232_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6216_ (.A1(_1812_),
    .A2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6217_ (.A1(_1137_),
    .A2(_2059_),
    .B(_2005_),
    .C(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6218_ (.A1(_1869_),
    .A2(_2229_),
    .B(_2235_),
    .C(_2008_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6219_ (.I(_1251_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6220_ (.I0(\as2650.stack[7][7] ),
    .I1(\as2650.stack[4][7] ),
    .I2(\as2650.stack[5][7] ),
    .I3(\as2650.stack[6][7] ),
    .S0(_0928_),
    .S1(_2237_),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_1457_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6222_ (.A1(_2199_),
    .A2(\as2650.stack[1][7] ),
    .B1(\as2650.stack[0][7] ),
    .B2(_1252_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6223_ (.I(_1919_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6224_ (.A1(_1209_),
    .A2(\as2650.stack[3][7] ),
    .B1(\as2650.stack[2][7] ),
    .B2(_2241_),
    .C(_2162_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6225_ (.A1(_2239_),
    .A2(_2240_),
    .B(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6226_ (.A1(_2159_),
    .A2(_2238_),
    .B(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6227_ (.A1(_1429_),
    .A2(_2210_),
    .B1(_2244_),
    .B2(_1927_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6228_ (.A1(_2217_),
    .A2(_2218_),
    .A3(_2236_),
    .B(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6229_ (.A1(_2210_),
    .A2(_2219_),
    .B1(_2246_),
    .B2(_2206_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6230_ (.A1(_2129_),
    .A2(_2247_),
    .B(_2127_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6231_ (.A1(_0972_),
    .A2(_1936_),
    .B(_2248_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6232_ (.I(_1735_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6233_ (.I(_1798_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6234_ (.A1(_0970_),
    .A2(_2209_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6235_ (.A1(_0974_),
    .A2(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6236_ (.A1(_2173_),
    .A2(_2212_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6237_ (.I(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6238_ (.A1(_0969_),
    .A2(_0538_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6239_ (.A1(_2176_),
    .A2(_2254_),
    .B(_2255_),
    .C(_2213_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6240_ (.A1(_2085_),
    .A2(_2090_),
    .A3(_2132_),
    .A4(_2254_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6241_ (.A1(\as2650.pc[8] ),
    .A2(_1185_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6242_ (.A1(_2256_),
    .A2(_2257_),
    .B(_2258_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6243_ (.A1(_2258_),
    .A2(_2256_),
    .A3(_2257_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6244_ (.A1(_2259_),
    .A2(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6245_ (.A1(_2211_),
    .A2(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6246_ (.A1(_1902_),
    .A2(_2252_),
    .B(_2262_),
    .C(_1572_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6247_ (.I(_0857_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6248_ (.A1(_2264_),
    .A2(_2261_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6249_ (.I(_0817_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6250_ (.A1(_1432_),
    .A2(_2252_),
    .B(_2265_),
    .C(_2266_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6251_ (.I(_3281_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6252_ (.A1(_1525_),
    .A2(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6253_ (.A1(_1915_),
    .A2(_2269_),
    .B(_1441_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6254_ (.A1(_1234_),
    .A2(_2221_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6255_ (.A1(_0975_),
    .A2(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6256_ (.A1(_0869_),
    .A2(_2267_),
    .A3(_2270_),
    .B1(_2220_),
    .B2(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6257_ (.I(\as2650.addr_buff[0] ),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6258_ (.I(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6259_ (.A1(net3),
    .A2(_3341_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6260_ (.A1(_1134_),
    .A2(_3341_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6261_ (.A1(_2232_),
    .A2(_2276_),
    .B(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_3280_),
    .A2(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6263_ (.A1(_2275_),
    .A2(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6264_ (.A1(\as2650.addr_buff[0] ),
    .A2(_1498_),
    .A3(_2278_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6265_ (.A1(_2280_),
    .A2(_2281_),
    .B(_2060_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6266_ (.A1(_1655_),
    .A2(_2273_),
    .B(_2282_),
    .C(_1940_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6267_ (.A1(\as2650.stack[7][8] ),
    .A2(_1465_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6268_ (.A1(_1972_),
    .A2(\as2650.stack[5][8] ),
    .B1(\as2650.stack[4][8] ),
    .B2(_0897_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6269_ (.A1(_1457_),
    .A2(_2285_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6270_ (.A1(\as2650.stack[6][8] ),
    .A2(_2195_),
    .B1(_1922_),
    .B2(_2284_),
    .C(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(_1457_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6272_ (.A1(_2112_),
    .A2(\as2650.stack[1][8] ),
    .B1(\as2650.stack[0][8] ),
    .B2(_2237_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6273_ (.A1(_2119_),
    .A2(\as2650.stack[3][8] ),
    .B1(\as2650.stack[2][8] ),
    .B2(_2241_),
    .C(_2162_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6274_ (.A1(_2288_),
    .A2(_2289_),
    .B(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6275_ (.A1(_2122_),
    .A2(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6276_ (.A1(_0855_),
    .A2(_2252_),
    .B1(_2287_),
    .B2(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6277_ (.A1(_2263_),
    .A2(_2283_),
    .B1(_2293_),
    .B2(_1850_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6278_ (.A1(_2172_),
    .A2(_2263_),
    .B(_2180_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6279_ (.A1(_2250_),
    .A2(_2294_),
    .B1(_2295_),
    .B2(_2252_),
    .C(_1981_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6280_ (.A1(_0976_),
    .A2(_1886_),
    .B(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6281_ (.A1(_2249_),
    .A2(_2297_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6282_ (.A1(_0974_),
    .A2(_2251_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6283_ (.A1(_1240_),
    .A2(_2298_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6284_ (.A1(_1240_),
    .A2(_2230_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6285_ (.A1(_0979_),
    .A2(_1186_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6286_ (.A1(_2300_),
    .A2(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6287_ (.A1(\as2650.pc[8] ),
    .A2(_2230_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6288_ (.A1(_2303_),
    .A2(_2259_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6289_ (.A1(_2302_),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6290_ (.A1(_2211_),
    .A2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6291_ (.A1(_1902_),
    .A2(_2299_),
    .B(_2306_),
    .C(_1572_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6292_ (.A1(_2264_),
    .A2(_2305_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6293_ (.A1(_2053_),
    .A2(_2299_),
    .B(_2308_),
    .C(_0818_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(_1529_),
    .A2(_2268_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6295_ (.A1(_1960_),
    .A2(_2310_),
    .B(_1441_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6296_ (.A1(_0974_),
    .A2(_0969_),
    .A3(_2221_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6297_ (.A1(_0979_),
    .A2(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6298_ (.A1(_0869_),
    .A2(_2309_),
    .A3(_2311_),
    .B1(_2220_),
    .B2(_2313_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6299_ (.A1(_1528_),
    .A2(_2281_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6300_ (.A1(_2060_),
    .A2(_2315_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6301_ (.A1(_1655_),
    .A2(_2314_),
    .B(_2316_),
    .C(_1940_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6302_ (.A1(_2112_),
    .A2(\as2650.stack[1][9] ),
    .B1(\as2650.stack[0][9] ),
    .B2(_2237_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6303_ (.A1(_2119_),
    .A2(\as2650.stack[3][9] ),
    .B1(\as2650.stack[2][9] ),
    .B2(_2241_),
    .C(_1468_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6304_ (.A1(_2239_),
    .A2(_2318_),
    .B(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6305_ (.A1(_2112_),
    .A2(\as2650.stack[5][9] ),
    .B1(\as2650.stack[4][9] ),
    .B2(_2237_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6306_ (.A1(\as2650.stack[7][9] ),
    .A2(_1455_),
    .B1(_2241_),
    .B2(\as2650.stack[6][9] ),
    .C(_2074_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6307_ (.A1(_2288_),
    .A2(_2321_),
    .B(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6308_ (.A1(_2122_),
    .A2(_2320_),
    .A3(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6309_ (.A1(_0855_),
    .A2(_2299_),
    .B(_2324_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6310_ (.A1(_2307_),
    .A2(_2317_),
    .B1(_2325_),
    .B2(_1850_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6311_ (.A1(_2172_),
    .A2(_2307_),
    .B(_1799_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6312_ (.A1(_2250_),
    .A2(_2326_),
    .B1(_2327_),
    .B2(_2299_),
    .C(_1981_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6313_ (.A1(_1241_),
    .A2(_1984_),
    .B(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6314_ (.A1(_2249_),
    .A2(_2329_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6315_ (.A1(_1240_),
    .A2(\as2650.pc[8] ),
    .A3(_2251_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6316_ (.A1(\as2650.pc[10] ),
    .A2(_2330_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6317_ (.A1(_0985_),
    .A2(_0538_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6318_ (.I(_2332_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6319_ (.A1(_2303_),
    .A2(_2300_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6320_ (.A1(_2259_),
    .A2(_2302_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6321_ (.A1(_2334_),
    .A2(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6322_ (.A1(_2333_),
    .A2(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6323_ (.A1(_1989_),
    .A2(_2331_),
    .B1(_2337_),
    .B2(_1994_),
    .C(_1753_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6324_ (.A1(_2172_),
    .A2(_2338_),
    .B(_2180_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6325_ (.A1(_1535_),
    .A2(_2268_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6326_ (.A1(_1998_),
    .A2(_2340_),
    .B(_0839_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6327_ (.A1(_2264_),
    .A2(_2331_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6328_ (.A1(_1663_),
    .A2(_2337_),
    .B(_2342_),
    .C(_2266_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6329_ (.A1(_0979_),
    .A2(_2312_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6330_ (.A1(_1243_),
    .A2(_2344_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6331_ (.A1(_1707_),
    .A2(_2341_),
    .A3(_2343_),
    .B1(_2220_),
    .B2(_2345_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6332_ (.A1(_2274_),
    .A2(_1528_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6333_ (.A1(_2279_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6334_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2348_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6335_ (.A1(_2006_),
    .A2(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6336_ (.A1(_1782_),
    .A2(_2346_),
    .B(_2350_),
    .C(_1779_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6337_ (.A1(_2199_),
    .A2(\as2650.stack[5][10] ),
    .B1(\as2650.stack[4][10] ),
    .B2(_1252_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6338_ (.A1(\as2650.stack[7][10] ),
    .A2(_2115_),
    .B1(_1920_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6339_ (.A1(_2239_),
    .A2(_2352_),
    .B(_2353_),
    .C(_2162_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6340_ (.A1(_2199_),
    .A2(\as2650.stack[1][10] ),
    .B1(\as2650.stack[0][10] ),
    .B2(_1252_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6341_ (.A1(_1209_),
    .A2(\as2650.stack[3][10] ),
    .B1(\as2650.stack[2][10] ),
    .B2(_1920_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6342_ (.A1(_2239_),
    .A2(_2355_),
    .B(_2356_),
    .C(_1969_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6343_ (.A1(_0855_),
    .A2(_2354_),
    .A3(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6344_ (.A1(_0825_),
    .A2(_2331_),
    .B(_2358_),
    .C(_2034_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6345_ (.A1(_2338_),
    .A2(_2351_),
    .B(_2359_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6346_ (.A1(_2331_),
    .A2(_2339_),
    .B1(_2360_),
    .B2(_2206_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6347_ (.I(_0883_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6348_ (.A1(_2129_),
    .A2(_2361_),
    .B(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6349_ (.A1(_0987_),
    .A2(_1936_),
    .B(_2363_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6350_ (.A1(_1411_),
    .A2(\as2650.stack[1][11] ),
    .B1(\as2650.stack[0][11] ),
    .B2(_0898_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6351_ (.A1(_0894_),
    .A2(\as2650.stack[3][11] ),
    .B1(\as2650.stack[2][11] ),
    .B2(_2195_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6352_ (.A1(_1458_),
    .A2(_2364_),
    .B(_2365_),
    .C(_2159_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6353_ (.A1(_0929_),
    .A2(\as2650.stack[5][11] ),
    .B1(\as2650.stack[4][11] ),
    .B2(_0898_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6354_ (.A1(\as2650.stack[7][11] ),
    .A2(_2115_),
    .B1(_2195_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6355_ (.A1(_1458_),
    .A2(_2367_),
    .B(_2368_),
    .C(_1469_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6356_ (.A1(_2366_),
    .A2(_2369_),
    .B(_0867_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(_0985_),
    .A2(_2330_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6358_ (.A1(_1246_),
    .A2(_2371_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6359_ (.I(_2372_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6360_ (.A1(_0825_),
    .A2(_2373_),
    .B(_2034_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6361_ (.A1(_0989_),
    .A2(_2230_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6362_ (.A1(\as2650.pc[10] ),
    .A2(_0539_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6363_ (.A1(_2333_),
    .A2(_2336_),
    .B(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6364_ (.A1(_2375_),
    .A2(_2377_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6365_ (.A1(_1900_),
    .A2(_2378_),
    .B1(_2373_),
    .B2(_1903_),
    .C(_1462_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6366_ (.I0(_2378_),
    .I1(_2372_),
    .S(_0832_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6367_ (.A1(_1131_),
    .A2(_1739_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6368_ (.A1(\as2650.addr_buff[3] ),
    .A2(_0624_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6369_ (.A1(_2266_),
    .A2(_2381_),
    .A3(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6370_ (.A1(_1810_),
    .A2(_2380_),
    .B(_2383_),
    .C(_0822_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6371_ (.A1(_1243_),
    .A2(_2344_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6372_ (.A1(_0989_),
    .A2(_2385_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6373_ (.A1(_1767_),
    .A2(_2372_),
    .B1(_2386_),
    .B2(_2009_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6374_ (.A1(_2384_),
    .A2(_2387_),
    .B(_1640_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6375_ (.I(\as2650.addr_buff[3] ),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6376_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6377_ (.A1(_2279_),
    .A2(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6378_ (.A1(_2389_),
    .A2(_2391_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6379_ (.A1(_1426_),
    .A2(_2373_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6380_ (.A1(_1761_),
    .A2(_2392_),
    .B1(_2393_),
    .B2(_2006_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6381_ (.A1(_1319_),
    .A2(_2388_),
    .A3(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6382_ (.A1(_2370_),
    .A2(_2374_),
    .B1(_2379_),
    .B2(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6383_ (.A1(_1800_),
    .A2(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6384_ (.A1(_1888_),
    .A2(_2373_),
    .B(_1889_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6385_ (.A1(_0990_),
    .A2(_1886_),
    .B1(_2397_),
    .B2(_2398_),
    .C(_1591_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6386_ (.A1(_1246_),
    .A2(_2371_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6387_ (.A1(_0993_),
    .A2(_2399_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6388_ (.I(_2400_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6389_ (.I(_1300_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6390_ (.A1(_1562_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6391_ (.A1(_2332_),
    .A2(_2375_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6392_ (.A1(_1246_),
    .A2(_0539_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6393_ (.A1(_2303_),
    .A2(_2300_),
    .A3(_2376_),
    .A4(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6394_ (.A1(_2335_),
    .A2(_2404_),
    .B(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6395_ (.A1(\as2650.pc[12] ),
    .A2(_0540_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6396_ (.A1(_2407_),
    .A2(_2408_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_1899_),
    .A2(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6398_ (.A1(_2403_),
    .A2(_2401_),
    .B(_2410_),
    .C(_1452_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6399_ (.A1(_1247_),
    .A2(_1243_),
    .A3(_2344_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6400_ (.A1(_1249_),
    .A2(_2412_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6401_ (.I(_2401_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6402_ (.A1(_1426_),
    .A2(_1893_),
    .A3(_2413_),
    .B1(_2414_),
    .B2(_1895_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6403_ (.A1(_2389_),
    .A2(_2279_),
    .A3(_2390_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6404_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2416_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6405_ (.A1(_2264_),
    .A2(_2400_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6406_ (.A1(_2053_),
    .A2(_2409_),
    .B(_2418_),
    .C(_1052_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(\as2650.addr_buff[4] ),
    .A2(_1945_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6408_ (.A1(_0378_),
    .A2(_1424_),
    .B(_1671_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6409_ (.A1(_2420_),
    .A2(_2421_),
    .B(_1639_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6410_ (.A1(_1517_),
    .A2(_2417_),
    .B1(_2419_),
    .B2(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6411_ (.A1(_1718_),
    .A2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6412_ (.A1(_2415_),
    .A2(_2424_),
    .B(_1765_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6413_ (.A1(_1212_),
    .A2(\as2650.stack[5][12] ),
    .B1(\as2650.stack[4][12] ),
    .B2(_2072_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6414_ (.A1(\as2650.stack[7][12] ),
    .A2(_1455_),
    .B1(_1974_),
    .B2(\as2650.stack[6][12] ),
    .C(_1968_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6415_ (.A1(_2288_),
    .A2(_2426_),
    .B(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6416_ (.A1(_1212_),
    .A2(\as2650.stack[1][12] ),
    .B1(\as2650.stack[0][12] ),
    .B2(_2072_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6417_ (.A1(_2119_),
    .A2(\as2650.stack[3][12] ),
    .B1(\as2650.stack[2][12] ),
    .B2(_1929_),
    .C(_1468_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6418_ (.A1(_2288_),
    .A2(_2429_),
    .B(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6419_ (.A1(_0824_),
    .A2(_2428_),
    .A3(_2431_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6420_ (.A1(_0867_),
    .A2(_2401_),
    .B(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6421_ (.A1(_2411_),
    .A2(_2425_),
    .B1(_2433_),
    .B2(_1453_),
    .C(_1939_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6422_ (.A1(_1888_),
    .A2(_2401_),
    .B(_2434_),
    .C(_1981_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6423_ (.A1(_0994_),
    .A2(_1886_),
    .B(_2435_),
    .C(_1695_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6424_ (.A1(_1081_),
    .A2(_0838_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6425_ (.A1(_2436_),
    .A2(_1593_),
    .B1(_1602_),
    .B2(_1606_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6426_ (.A1(_0655_),
    .A2(_0637_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6427_ (.A1(_3206_),
    .A2(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6428_ (.A1(_3237_),
    .A2(_3240_),
    .B(_2439_),
    .C(_3350_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6429_ (.A1(_0679_),
    .A2(_1010_),
    .B(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6430_ (.A1(_0648_),
    .A2(_2441_),
    .B(_1030_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6431_ (.A1(_3236_),
    .A2(_3240_),
    .B1(_3281_),
    .B2(_3276_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6432_ (.A1(_1437_),
    .A2(_2443_),
    .B(_3304_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6433_ (.A1(_1080_),
    .A2(_1006_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6434_ (.A1(_1025_),
    .A2(_3266_),
    .A3(_0655_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6435_ (.A1(_1063_),
    .A2(_2445_),
    .B1(_2446_),
    .B2(_1501_),
    .C(_1613_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6436_ (.A1(_1055_),
    .A2(_1058_),
    .A3(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6437_ (.A1(_3202_),
    .A2(_3310_),
    .A3(_1008_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6438_ (.A1(_3156_),
    .A2(_1043_),
    .B(_1686_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6439_ (.A1(_1869_),
    .A2(_1047_),
    .A3(_2449_),
    .A4(_2450_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6440_ (.A1(_1034_),
    .A2(_1021_),
    .A3(_1038_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6441_ (.A1(_2444_),
    .A2(_2448_),
    .A3(_2451_),
    .A4(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6442_ (.A1(_2437_),
    .A2(_2442_),
    .A3(_2453_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_2454_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6444_ (.A1(_3317_),
    .A2(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6445_ (.I(_1004_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6446_ (.I(_1682_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6447_ (.A1(_2458_),
    .A2(_3303_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6448_ (.A1(_1827_),
    .A2(_3391_),
    .B(_2459_),
    .C(_1768_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6449_ (.A1(_1760_),
    .A2(_3446_),
    .B(_2457_),
    .C(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6450_ (.I(_3438_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6451_ (.I(_1145_),
    .Z(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6452_ (.I(_1046_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6453_ (.I(_1114_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6454_ (.A1(_0844_),
    .A2(_1099_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6456_ (.A1(_3432_),
    .A2(_2467_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6457_ (.I(_0846_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6458_ (.A1(\as2650.psu[0] ),
    .A2(_2469_),
    .B(_1114_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6459_ (.I(_0806_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6460_ (.A1(_2465_),
    .A2(_3348_),
    .B1(_2468_),
    .B2(_2470_),
    .C(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6461_ (.A1(_1096_),
    .A2(_3362_),
    .B(_1158_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6462_ (.A1(_1128_),
    .A2(_1138_),
    .B1(_2472_),
    .B2(_2473_),
    .C(_1504_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6463_ (.A1(_2462_),
    .A2(_2463_),
    .B1(_2464_),
    .B2(_3370_),
    .C(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6464_ (.I(_2454_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6465_ (.A1(_2461_),
    .A2(_2475_),
    .A3(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6466_ (.A1(_1650_),
    .A2(_2456_),
    .A3(_2477_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6467_ (.I(_2454_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6468_ (.I(_1082_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6469_ (.A1(_2458_),
    .A2(_3527_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6470_ (.A1(_1855_),
    .A2(_3492_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6471_ (.A1(_1436_),
    .A2(_2480_),
    .A3(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6472_ (.A1(_1741_),
    .A2(_3484_),
    .B(_2479_),
    .C(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6473_ (.A1(_1064_),
    .A2(_0847_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6474_ (.A1(\as2650.psu[1] ),
    .A2(_2466_),
    .B(_1097_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6475_ (.A1(_1652_),
    .A2(_2462_),
    .B1(_2484_),
    .B2(_2485_),
    .C(_1095_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6476_ (.A1(_0806_),
    .A2(_0726_),
    .B(_3223_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6477_ (.A1(_1129_),
    .A2(_1123_),
    .B1(_2486_),
    .B2(_2487_),
    .C(_1412_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6478_ (.A1(_1413_),
    .A2(_3514_),
    .B(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6479_ (.A1(_1118_),
    .A2(_1854_),
    .B1(_2489_),
    .B2(_1204_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6480_ (.A1(_2478_),
    .A2(_2483_),
    .A3(_2490_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6481_ (.A1(_3494_),
    .A2(_2476_),
    .B(_2491_),
    .C(_1695_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6482_ (.A1(_1713_),
    .A2(_2455_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6483_ (.I(_1436_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6484_ (.I(_1682_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6485_ (.A1(_2494_),
    .A2(_3545_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6486_ (.A1(_1856_),
    .A2(_3552_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6487_ (.A1(_2493_),
    .A2(_2495_),
    .A3(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6488_ (.I(_1154_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6489_ (.A1(_0751_),
    .A2(_0278_),
    .B(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6490_ (.A1(\as2650.overflow ),
    .A2(_2466_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6491_ (.A1(_1183_),
    .A2(_2467_),
    .B(_2500_),
    .C(_1097_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6492_ (.A1(_1098_),
    .A2(_1118_),
    .B(_2501_),
    .C(_1121_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6493_ (.A1(_1096_),
    .A2(_0741_),
    .B(_2502_),
    .C(_1158_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6494_ (.A1(_1534_),
    .A2(_1123_),
    .B(_1633_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6495_ (.A1(_0321_),
    .A2(_1554_),
    .B1(_2503_),
    .B2(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6496_ (.A1(_3567_),
    .A2(_2464_),
    .B(_2478_),
    .C(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6497_ (.A1(_2497_),
    .A2(_2499_),
    .B(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6498_ (.A1(_1650_),
    .A2(_2492_),
    .A3(_2507_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6499_ (.A1(_0725_),
    .A2(_2455_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6500_ (.I(_2454_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6501_ (.I(_1425_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6502_ (.A1(_1683_),
    .A2(_0313_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6503_ (.A1(_1827_),
    .A2(_0349_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6504_ (.A1(_2510_),
    .A2(_2511_),
    .A3(_2512_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6505_ (.A1(_1741_),
    .A2(_0307_),
    .B(_2479_),
    .C(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6506_ (.A1(_0334_),
    .A2(_1665_),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6507_ (.I(_1095_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6508_ (.A1(_3326_),
    .A2(_0847_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6509_ (.A1(\as2650.psu[3] ),
    .A2(_2467_),
    .B(_1652_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6510_ (.A1(_1098_),
    .A2(_0726_),
    .B1(_2517_),
    .B2(_2518_),
    .C(_1121_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6511_ (.A1(_2516_),
    .A2(_0482_),
    .B(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6512_ (.A1(_1159_),
    .A2(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6513_ (.I(_1123_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6514_ (.A1(_1537_),
    .A2(_2522_),
    .B(_1633_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6515_ (.A1(_0365_),
    .A2(_1854_),
    .B1(_2521_),
    .B2(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6516_ (.A1(_2509_),
    .A2(_2514_),
    .A3(_2515_),
    .A4(_2524_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6517_ (.A1(_1650_),
    .A2(_2508_),
    .A3(_2525_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6518_ (.A1(_0363_),
    .A2(_2509_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(_2494_),
    .A2(_0362_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(_1856_),
    .A2(_0391_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6521_ (.A1(_2493_),
    .A2(_2527_),
    .A3(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6522_ (.A1(_0751_),
    .A2(_0423_),
    .B(_2457_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6523_ (.A1(\as2650.psu[4] ),
    .A2(_2469_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6524_ (.A1(_3335_),
    .A2(_0848_),
    .B(_2531_),
    .C(_1653_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6525_ (.A1(_1653_),
    .A2(_0365_),
    .B(_2532_),
    .C(_2516_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6526_ (.A1(_2516_),
    .A2(_0772_),
    .B(_2533_),
    .C(_1159_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6527_ (.A1(_1541_),
    .A2(_2522_),
    .B(_1634_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6528_ (.A1(_0472_),
    .A2(_2463_),
    .B1(_1665_),
    .B2(_0381_),
    .C(_2478_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6529_ (.A1(_2529_),
    .A2(_2530_),
    .B1(_2534_),
    .B2(_2535_),
    .C(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6530_ (.A1(_1150_),
    .A2(_2526_),
    .A3(_2537_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6531_ (.A1(_0471_),
    .A2(_2509_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6532_ (.A1(_2471_),
    .A2(_0586_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6533_ (.A1(_2465_),
    .A2(_0482_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6534_ (.A1(_2539_),
    .A2(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6535_ (.A1(\as2650.psu[5] ),
    .A2(_2467_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6536_ (.A1(\as2650.psl[5] ),
    .A2(_0848_),
    .B(_2542_),
    .C(_0808_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6537_ (.A1(_1159_),
    .A2(_2541_),
    .A3(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6538_ (.A1(_1544_),
    .A2(_2522_),
    .B(_1634_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6539_ (.A1(_0772_),
    .A2(_2463_),
    .B1(_2464_),
    .B2(_0488_),
    .C(_2478_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6540_ (.A1(_1683_),
    .A2(_0467_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6541_ (.A1(_2494_),
    .A2(_0470_),
    .B(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6542_ (.A1(_2510_),
    .A2(_0453_),
    .B(_1083_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6543_ (.A1(_2493_),
    .A2(_2548_),
    .B(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6544_ (.A1(_2544_),
    .A2(_2545_),
    .B(_2546_),
    .C(_2550_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6545_ (.A1(_1150_),
    .A2(_2538_),
    .A3(_2551_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6546_ (.A1(_1728_),
    .A2(_2455_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6547_ (.A1(_1683_),
    .A2(_0535_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_1855_),
    .A2(_0549_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6549_ (.A1(_2510_),
    .A2(_2553_),
    .A3(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6550_ (.A1(_1741_),
    .A2(_0528_),
    .B(_2479_),
    .C(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6551_ (.A1(net27),
    .A2(_0847_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6552_ (.A1(_0997_),
    .A2(_2469_),
    .B(_2557_),
    .C(_1652_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6553_ (.A1(_1098_),
    .A2(_0448_),
    .B(_2558_),
    .C(_1096_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6554_ (.A1(_2516_),
    .A2(_1141_),
    .B(_2559_),
    .C(_1138_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6555_ (.A1(_1546_),
    .A2(_2522_),
    .B(_1633_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6556_ (.A1(_0586_),
    .A2(_1854_),
    .B1(_2560_),
    .B2(_2561_),
    .C(_2476_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6557_ (.A1(_0537_),
    .A2(_2464_),
    .B(_2556_),
    .C(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6558_ (.A1(_1151_),
    .A2(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6559_ (.A1(_2552_),
    .A2(_2564_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6560_ (.A1(_0585_),
    .A2(_2509_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6561_ (.A1(_2494_),
    .A2(_0583_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6562_ (.A1(_1856_),
    .A2(_0600_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6563_ (.A1(_2493_),
    .A2(_2566_),
    .A3(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6564_ (.A1(_2510_),
    .A2(_0577_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6565_ (.A1(_2498_),
    .A2(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6566_ (.A1(_1160_),
    .A2(_2469_),
    .B(_0808_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6567_ (.A1(_1182_),
    .A2(_0848_),
    .B(_2571_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6568_ (.A1(_1157_),
    .A2(_1138_),
    .B1(_1202_),
    .B2(_2572_),
    .C(_1504_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6569_ (.A1(_1141_),
    .A2(_2463_),
    .B1(_1665_),
    .B2(_0591_),
    .C(_2573_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6570_ (.A1(_2568_),
    .A2(_2570_),
    .B(_2574_),
    .C(_2476_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6571_ (.A1(_1150_),
    .A2(_2565_),
    .A3(_2575_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6572_ (.A1(_0895_),
    .A2(_0899_),
    .A3(_1214_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6573_ (.I(_2576_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6574_ (.I(_2577_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6575_ (.I(_2576_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6576_ (.A1(\as2650.stack[7][0] ),
    .A2(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6577_ (.A1(_0891_),
    .A2(_2578_),
    .B(_2580_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6578_ (.A1(\as2650.stack[7][1] ),
    .A2(_2579_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6579_ (.A1(_0938_),
    .A2(_2578_),
    .B(_2581_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6580_ (.A1(\as2650.stack[7][2] ),
    .A2(_2579_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6581_ (.A1(_0944_),
    .A2(_2578_),
    .B(_2582_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6582_ (.A1(\as2650.stack[7][3] ),
    .A2(_2579_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6583_ (.A1(_0950_),
    .A2(_2578_),
    .B(_2583_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6584_ (.I(_2577_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6585_ (.I(_2576_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6586_ (.A1(\as2650.stack[7][4] ),
    .A2(_2585_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6587_ (.A1(_0954_),
    .A2(_2584_),
    .B(_2586_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6588_ (.A1(\as2650.stack[7][5] ),
    .A2(_2585_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6589_ (.A1(_0961_),
    .A2(_2584_),
    .B(_2587_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6590_ (.A1(\as2650.stack[7][6] ),
    .A2(_2585_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6591_ (.A1(_0966_),
    .A2(_2584_),
    .B(_2588_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(\as2650.stack[7][7] ),
    .A2(_2585_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6593_ (.A1(_0971_),
    .A2(_2584_),
    .B(_2589_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6594_ (.I0(_1237_),
    .I1(\as2650.stack[7][8] ),
    .S(_2577_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(_2590_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6596_ (.I(_2577_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6597_ (.I(_2576_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6598_ (.A1(\as2650.stack[7][9] ),
    .A2(_2592_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6599_ (.A1(_0980_),
    .A2(_2591_),
    .B(_2593_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(\as2650.stack[7][10] ),
    .A2(_2592_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6601_ (.A1(_0986_),
    .A2(_2591_),
    .B(_2594_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6602_ (.A1(\as2650.stack[7][11] ),
    .A2(_2592_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6603_ (.A1(_0990_),
    .A2(_2591_),
    .B(_2595_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6604_ (.A1(\as2650.stack[7][12] ),
    .A2(_2592_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6605_ (.A1(_0994_),
    .A2(_2591_),
    .B(_2596_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(net28),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6607_ (.A1(_0901_),
    .A2(_1517_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6608_ (.A1(_1514_),
    .A2(_2598_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6609_ (.A1(_1420_),
    .A2(_1551_),
    .A3(_1046_),
    .A4(_1578_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6610_ (.A1(_1034_),
    .A2(_2599_),
    .B(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6611_ (.A1(_1587_),
    .A2(_1617_),
    .A3(_1685_),
    .A4(_1874_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6612_ (.A1(_1503_),
    .A2(_1599_),
    .A3(_1882_),
    .A4(_2602_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6613_ (.A1(_1419_),
    .A2(_2601_),
    .B(_2603_),
    .C(_1597_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6614_ (.A1(_1631_),
    .A2(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(_2605_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_2606_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6617_ (.I(_1579_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6618_ (.I(_1742_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6619_ (.A1(_2609_),
    .A2(_1898_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6620_ (.I(_1493_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(_2611_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6622_ (.A1(_1420_),
    .A2(_3236_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6623_ (.A1(_3391_),
    .A2(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6624_ (.A1(_1487_),
    .A2(_2614_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6625_ (.A1(_3267_),
    .A2(_3303_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6626_ (.I(_1495_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6627_ (.A1(_1907_),
    .A2(_2616_),
    .B(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6628_ (.A1(_1907_),
    .A2(_2616_),
    .B(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6629_ (.A1(_2458_),
    .A2(_2615_),
    .B(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6630_ (.A1(_2597_),
    .A2(_2612_),
    .B1(_2620_),
    .B2(_1600_),
    .C(_1154_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6631_ (.A1(_1439_),
    .A2(_0868_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6632_ (.I(_2622_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6633_ (.A1(_2597_),
    .A2(_1425_),
    .B(_1909_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6634_ (.A1(_0900_),
    .A2(_1299_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6635_ (.I(_2625_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6636_ (.A1(_2402_),
    .A2(_1898_),
    .B1(_2624_),
    .B2(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6637_ (.A1(_2266_),
    .A2(_1427_),
    .B(_2622_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6638_ (.A1(_2623_),
    .A2(_2627_),
    .B1(_2628_),
    .B2(_0890_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6639_ (.A1(_2610_),
    .A2(_2621_),
    .B1(_2629_),
    .B2(_1204_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6640_ (.A1(_1145_),
    .A2(_1645_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6641_ (.A1(_1208_),
    .A2(_2631_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6642_ (.A1(_2608_),
    .A2(_2630_),
    .B(_2632_),
    .C(_2606_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6643_ (.A1(_2597_),
    .A2(_2607_),
    .B(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6644_ (.A1(_2249_),
    .A2(_2634_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(_2606_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6646_ (.A1(_1554_),
    .A2(_1579_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(_2636_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6648_ (.I(_1787_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6649_ (.A1(net52),
    .A2(net28),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_3309_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6651_ (.I(_2640_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6652_ (.A1(_3371_),
    .A2(_3302_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6653_ (.A1(_1171_),
    .A2(_3486_),
    .A3(_3524_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6654_ (.A1(_2642_),
    .A2(_2643_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6655_ (.A1(_3507_),
    .A2(_2640_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6656_ (.A1(_0317_),
    .A2(_1605_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6657_ (.A1(_1746_),
    .A2(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(_2647_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6659_ (.A1(_2641_),
    .A2(_2644_),
    .B(_2645_),
    .C(_2648_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6660_ (.A1(_3371_),
    .A2(_3390_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6661_ (.A1(_1171_),
    .A2(_3486_),
    .A3(_3489_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6662_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3235_),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6663_ (.I(_2652_),
    .Z(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6664_ (.A1(_2650_),
    .A2(_2651_),
    .B(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6665_ (.A1(_2650_),
    .A2(_2651_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6666_ (.A1(_1173_),
    .A2(_2613_),
    .B(_2655_),
    .C(_1826_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6667_ (.A1(_2649_),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6668_ (.A1(_0317_),
    .A2(_1488_),
    .A3(_1489_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6669_ (.A1(_1842_),
    .A2(_2658_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6670_ (.A1(_2612_),
    .A2(_2639_),
    .B1(_2657_),
    .B2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6671_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6672_ (.A1(_2661_),
    .A2(_1950_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6673_ (.A1(_2661_),
    .A2(_1950_),
    .B(_1788_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6674_ (.A1(_2638_),
    .A2(_2660_),
    .B1(_2662_),
    .B2(_2663_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6675_ (.I(_2628_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_1300_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6677_ (.I(_1498_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6678_ (.A1(_1768_),
    .A2(_2639_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6679_ (.A1(_1129_),
    .A2(_2667_),
    .B(_2668_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6680_ (.A1(_2666_),
    .A2(_1951_),
    .B1(_2669_),
    .B2(_2626_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6681_ (.A1(_1219_),
    .A2(_2665_),
    .B1(_2670_),
    .B2(_2623_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6682_ (.A1(_1084_),
    .A2(_2664_),
    .B1(_2671_),
    .B2(_1094_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6683_ (.A1(_1219_),
    .A2(_2637_),
    .B1(_2672_),
    .B2(_2608_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6684_ (.I(_2605_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6685_ (.A1(net29),
    .A2(_2674_),
    .B(_2362_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6686_ (.A1(_2635_),
    .A2(_2673_),
    .B(_2675_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6687_ (.I(net30),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6688_ (.I(_2605_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_2677_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6690_ (.A1(_1172_),
    .A2(_3525_),
    .A3(_3526_),
    .B1(_2642_),
    .B2(_2643_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6691_ (.A1(_3570_),
    .A2(_3545_),
    .A3(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6692_ (.A1(_2641_),
    .A2(_2680_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_3267_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6694_ (.A1(_1130_),
    .A2(_2682_),
    .B(_2648_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6695_ (.I(_2653_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6696_ (.A1(_1172_),
    .A2(_3490_),
    .A3(_3491_),
    .B1(_2650_),
    .B2(_2651_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6697_ (.A1(_3570_),
    .A2(_3552_),
    .A3(_2685_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6698_ (.I(_2652_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6699_ (.A1(_1534_),
    .A2(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6700_ (.A1(_2684_),
    .A2(_2686_),
    .B(_2688_),
    .C(_1826_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6701_ (.A1(_2681_),
    .A2(_2683_),
    .B(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6702_ (.A1(net52),
    .A2(_2597_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6703_ (.A1(_2676_),
    .A2(_2691_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_2611_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6705_ (.A1(_1991_),
    .A2(_2662_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6706_ (.A1(_1990_),
    .A2(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6707_ (.A1(_1600_),
    .A2(_2690_),
    .B1(_2692_),
    .B2(_2693_),
    .C1(_2695_),
    .C2(_1847_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6708_ (.A1(_2498_),
    .A2(_1579_),
    .A3(_2696_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6709_ (.I(_2631_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6710_ (.A1(_1461_),
    .A2(_2018_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6711_ (.A1(_1568_),
    .A2(_2666_),
    .B(_2699_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6712_ (.A1(_1801_),
    .A2(_2692_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6713_ (.A1(_2015_),
    .A2(_2701_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6714_ (.A1(_1664_),
    .A2(_2012_),
    .B1(_2702_),
    .B2(_1672_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6715_ (.A1(_0943_),
    .A2(_2700_),
    .B1(_2703_),
    .B2(_2699_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6716_ (.I(_2677_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6717_ (.A1(_0942_),
    .A2(_2698_),
    .B1(_2704_),
    .B2(_1800_),
    .C(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6718_ (.A1(_2676_),
    .A2(_2678_),
    .B1(_2697_),
    .B2(_2706_),
    .C(_1591_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6719_ (.I(net31),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6720_ (.A1(_1990_),
    .A2(_2694_),
    .B(_2044_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6721_ (.A1(_2042_),
    .A2(_2708_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6722_ (.A1(net30),
    .A2(net52),
    .A3(net28),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6723_ (.A1(_2707_),
    .A2(_2710_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6724_ (.I(_0336_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6725_ (.A1(_3539_),
    .A2(_3542_),
    .A3(_3544_),
    .B(_1533_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6726_ (.A1(_1533_),
    .A2(_3539_),
    .A3(_3542_),
    .A4(_3544_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6727_ (.A1(_2679_),
    .A2(_2713_),
    .B(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6728_ (.A1(_2712_),
    .A2(_0313_),
    .A3(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6729_ (.A1(_3310_),
    .A2(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6730_ (.A1(_1131_),
    .A2(_3310_),
    .B(_2617_),
    .C(_2717_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6731_ (.A1(_3547_),
    .A2(_3549_),
    .A3(_3551_),
    .B(_1533_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6732_ (.A1(_1532_),
    .A2(_3547_),
    .A3(_3549_),
    .A4(_3551_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6733_ (.A1(_2685_),
    .A2(_2719_),
    .B(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6734_ (.A1(_0337_),
    .A2(_0349_),
    .A3(_2721_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6735_ (.A1(_2653_),
    .A2(_2722_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6736_ (.A1(_1131_),
    .A2(_2653_),
    .B(_2723_),
    .C(_1492_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6737_ (.A1(_2718_),
    .A2(_2724_),
    .B(_2659_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6738_ (.A1(_1605_),
    .A2(_2711_),
    .B(_2725_),
    .C(_1787_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6739_ (.A1(_1788_),
    .A2(_2709_),
    .B(_2726_),
    .C(_1083_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6740_ (.A1(_1739_),
    .A2(_2711_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6741_ (.A1(_1174_),
    .A2(_1801_),
    .B(_2728_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6742_ (.A1(_1040_),
    .A2(_2402_),
    .A3(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6743_ (.A1(_1414_),
    .A2(_2402_),
    .B(_0839_),
    .C(_1222_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6744_ (.A1(_1833_),
    .A2(_2047_),
    .A3(_2730_),
    .A4(_2731_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6745_ (.A1(_1222_),
    .A2(_1634_),
    .B(_2727_),
    .C(_2732_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6746_ (.A1(_0949_),
    .A2(_2631_),
    .B1(_2733_),
    .B2(_1646_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6747_ (.A1(_2705_),
    .A2(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6748_ (.I(_1472_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6749_ (.A1(_2707_),
    .A2(_2678_),
    .B(_2735_),
    .C(_2736_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6750_ (.A1(_2087_),
    .A2(_2708_),
    .B(_2088_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6751_ (.A1(_2086_),
    .A2(_2737_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6752_ (.I(net32),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6753_ (.A1(_2707_),
    .A2(_2710_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6754_ (.A1(_2739_),
    .A2(_2740_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6755_ (.A1(_2712_),
    .A2(_0348_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6756_ (.A1(_0336_),
    .A2(_0348_),
    .B1(_2685_),
    .B2(_2719_),
    .C(_2720_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6757_ (.A1(_2742_),
    .A2(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6758_ (.A1(_1540_),
    .A2(_0391_),
    .A3(_2744_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6759_ (.A1(_2613_),
    .A2(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6760_ (.A1(_1540_),
    .A2(_2684_),
    .B(_0318_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6761_ (.A1(_1184_),
    .A2(_0361_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6762_ (.A1(_2712_),
    .A2(_0312_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6763_ (.A1(_2712_),
    .A2(_0312_),
    .B1(_2679_),
    .B2(_2713_),
    .C(_2714_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6764_ (.A1(_2749_),
    .A2(_2750_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6765_ (.A1(_2748_),
    .A2(_2751_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6766_ (.A1(_0378_),
    .A2(_3267_),
    .B(_2647_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6767_ (.A1(_2682_),
    .A2(_2752_),
    .B(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6768_ (.A1(_2746_),
    .A2(_2747_),
    .B(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6769_ (.A1(_2658_),
    .A2(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6770_ (.A1(_1857_),
    .A2(_2738_),
    .B1(_2741_),
    .B2(_2693_),
    .C(_2756_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6771_ (.A1(_2268_),
    .A2(_2741_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6772_ (.A1(_1540_),
    .A2(_1499_),
    .B(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6773_ (.A1(_2625_),
    .A2(_2759_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6774_ (.A1(_1940_),
    .A2(_2091_),
    .B(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6775_ (.A1(_1226_),
    .A2(_2700_),
    .B1(_2761_),
    .B2(_2699_),
    .C(_1755_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6776_ (.A1(_2498_),
    .A2(_2757_),
    .B(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6777_ (.A1(_1226_),
    .A2(_2698_),
    .B1(_2763_),
    .B2(_1690_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6778_ (.A1(_2739_),
    .A2(_2674_),
    .B(_2362_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6779_ (.A1(_2635_),
    .A2(_2764_),
    .B(_2765_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6780_ (.A1(_2086_),
    .A2(_2737_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6781_ (.A1(_2134_),
    .A2(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6782_ (.A1(_2133_),
    .A2(_2767_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6783_ (.I(_1606_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6784_ (.A1(_0872_),
    .A2(_2684_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6785_ (.A1(_0388_),
    .A2(_0390_),
    .B(_0375_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6786_ (.A1(_0376_),
    .A2(_0388_),
    .A3(_0390_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6787_ (.A1(_2742_),
    .A2(_2771_),
    .A3(_2743_),
    .B(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6788_ (.A1(_0871_),
    .A2(_0470_),
    .A3(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6789_ (.A1(_2613_),
    .A2(_2774_),
    .B(_1682_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6790_ (.A1(_0376_),
    .A2(_0362_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6791_ (.A1(_2749_),
    .A2(_2748_),
    .A3(_2750_),
    .B(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6792_ (.A1(_0760_),
    .A2(_0467_),
    .A3(_2777_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6793_ (.A1(_1544_),
    .A2(_2682_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6794_ (.A1(_2682_),
    .A2(_2778_),
    .B(_2779_),
    .C(_2617_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6795_ (.A1(_2770_),
    .A2(_2775_),
    .B(_2780_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6796_ (.A1(_2739_),
    .A2(_2740_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6797_ (.A1(net51),
    .A2(_2782_),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6798_ (.A1(_2611_),
    .A2(_2783_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6799_ (.A1(_2769_),
    .A2(_2781_),
    .B(_2784_),
    .C(_2638_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6800_ (.A1(_1821_),
    .A2(_2768_),
    .B(_2785_),
    .C(_1084_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(_2628_),
    .Z(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6802_ (.A1(_0872_),
    .A2(_1768_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6803_ (.A1(_2139_),
    .A2(_2783_),
    .B(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6804_ (.I(_1443_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6805_ (.A1(_1230_),
    .A2(_2787_),
    .B1(_2789_),
    .B2(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6806_ (.A1(_1900_),
    .A2(_2136_),
    .B(_2791_),
    .C(_2250_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6807_ (.A1(_1230_),
    .A2(_2637_),
    .B1(_2786_),
    .B2(_2608_),
    .C(_2792_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6808_ (.I(_2605_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6809_ (.A1(net33),
    .A2(_2794_),
    .B(_2362_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6810_ (.A1(_2635_),
    .A2(_2793_),
    .B(_2795_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6811_ (.A1(net51),
    .A2(_2739_),
    .A3(_2740_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6812_ (.A1(net34),
    .A2(_2796_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6813_ (.A1(_2693_),
    .A2(_2797_),
    .B(_1847_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6814_ (.I(_0489_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6815_ (.A1(_0454_),
    .A2(_0373_),
    .B1(_0460_),
    .B2(_0456_),
    .C(_0465_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6816_ (.A1(_2799_),
    .A2(_2800_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6817_ (.A1(_2799_),
    .A2(_2800_),
    .Z(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6818_ (.A1(_2777_),
    .A2(_2801_),
    .B(_2802_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6819_ (.A1(_1164_),
    .A2(_0535_),
    .A3(_2803_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6820_ (.A1(_2641_),
    .A2(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6821_ (.A1(_1126_),
    .A2(_2641_),
    .B(_2617_),
    .C(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6822_ (.A1(_1187_),
    .A2(_0548_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6823_ (.A1(_2799_),
    .A2(_0469_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6824_ (.A1(_2799_),
    .A2(_0469_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6825_ (.A1(_2808_),
    .A2(_2773_),
    .B(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6826_ (.A1(_2807_),
    .A2(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6827_ (.A1(_2807_),
    .A2(_2810_),
    .B(_2687_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6828_ (.A1(_1126_),
    .A2(_2684_),
    .B1(_2811_),
    .B2(_2812_),
    .C(_2458_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6829_ (.I(_2659_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6830_ (.A1(_2806_),
    .A2(_2813_),
    .B(_2814_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6831_ (.A1(_2133_),
    .A2(_2766_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6832_ (.A1(_2175_),
    .A2(_2816_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6833_ (.A1(_2173_),
    .A2(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6834_ (.A1(_2798_),
    .A2(_2815_),
    .B1(_2818_),
    .B2(_1857_),
    .C(_2457_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6835_ (.A1(_2667_),
    .A2(_2797_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6836_ (.A1(_1126_),
    .A2(_2139_),
    .B(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6837_ (.A1(_2666_),
    .A2(_2178_),
    .B1(_2821_),
    .B2(_2626_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6838_ (.A1(_1232_),
    .A2(_2665_),
    .B1(_2822_),
    .B2(_2623_),
    .C(_1582_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6839_ (.A1(_2819_),
    .A2(_2823_),
    .B(_1647_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6840_ (.A1(_1232_),
    .A2(_2637_),
    .B(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6841_ (.I(_0883_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6842_ (.A1(net34),
    .A2(_2794_),
    .B(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6843_ (.A1(_2635_),
    .A2(_2825_),
    .B(_2827_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6844_ (.I(net35),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6845_ (.A1(_0964_),
    .A2(_1109_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6846_ (.A1(_2829_),
    .A2(_2817_),
    .B(_2213_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6847_ (.A1(_2212_),
    .A2(_2830_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6848_ (.A1(net34),
    .A2(net51),
    .A3(net32),
    .A4(_2740_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6849_ (.A1(net35),
    .A2(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6850_ (.I(net3),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6851_ (.A1(_0540_),
    .A2(_0534_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6852_ (.A1(_1164_),
    .A2(_0534_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6853_ (.A1(_2835_),
    .A2(_2803_),
    .B(_2836_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6854_ (.A1(_2834_),
    .A2(_0582_),
    .A3(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6855_ (.A1(_1136_),
    .A2(_2640_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6856_ (.A1(_2640_),
    .A2(_2838_),
    .B(_2839_),
    .C(_2647_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6857_ (.A1(_1164_),
    .A2(_0549_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6858_ (.A1(_2807_),
    .A2(_2810_),
    .B(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6859_ (.A1(_2834_),
    .A2(_0599_),
    .A3(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6860_ (.A1(_1136_),
    .A2(_2687_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6861_ (.A1(_2687_),
    .A2(_2843_),
    .B(_2844_),
    .C(_1826_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6862_ (.A1(_2840_),
    .A2(_2845_),
    .B(_2769_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6863_ (.A1(_2612_),
    .A2(_2833_),
    .B(_2846_),
    .C(_1742_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6864_ (.A1(_2609_),
    .A2(_2831_),
    .B(_2847_),
    .C(_1154_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6865_ (.A1(_1760_),
    .A2(_2833_),
    .B(_2224_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6866_ (.A1(_1235_),
    .A2(_2787_),
    .B1(_2849_),
    .B2(_2790_),
    .C(_2217_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6867_ (.A1(_1235_),
    .A2(_2636_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6868_ (.A1(_1646_),
    .A2(_2848_),
    .B1(_2850_),
    .B2(_2250_),
    .C(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6869_ (.A1(_2705_),
    .A2(_2852_),
    .B(_2826_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6870_ (.A1(_2828_),
    .A2(_2678_),
    .B(_2853_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6871_ (.A1(_2254_),
    .A2(_2817_),
    .B(_2213_),
    .C(_2255_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6872_ (.A1(_2258_),
    .A2(_2854_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6873_ (.A1(_2258_),
    .A2(_2854_),
    .B(_2609_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6874_ (.A1(_0588_),
    .A2(_0582_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6875_ (.A1(_2835_),
    .A2(_2803_),
    .B(_2857_),
    .C(_2836_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6876_ (.A1(_2834_),
    .A2(_0583_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6877_ (.A1(_3309_),
    .A2(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6878_ (.A1(_2274_),
    .A2(_2858_),
    .A3(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6879_ (.A1(_2858_),
    .A2(_2860_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6880_ (.A1(_2275_),
    .A2(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6881_ (.A1(_2861_),
    .A2(_2863_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6882_ (.A1(_2834_),
    .A2(_0599_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6883_ (.A1(_2807_),
    .A2(_2810_),
    .B(_2865_),
    .C(_2841_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6884_ (.A1(_1135_),
    .A2(_0600_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6885_ (.A1(_2652_),
    .A2(_2867_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6886_ (.A1(_2274_),
    .A2(_2866_),
    .A3(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6887_ (.A1(_2866_),
    .A2(_2868_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6888_ (.A1(_2275_),
    .A2(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6889_ (.A1(_2869_),
    .A2(_2871_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6890_ (.A1(_2648_),
    .A2(_2864_),
    .B1(_2872_),
    .B2(_1855_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6891_ (.A1(_2828_),
    .A2(_2832_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6892_ (.A1(net50),
    .A2(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6893_ (.A1(_2611_),
    .A2(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6894_ (.A1(_2769_),
    .A2(_2873_),
    .B(_2876_),
    .C(_2638_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6895_ (.A1(_2855_),
    .A2(_2856_),
    .B(_1084_),
    .C(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6896_ (.A1(_2667_),
    .A2(_2875_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6897_ (.A1(_1525_),
    .A2(_0751_),
    .B(_2879_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6898_ (.A1(_1664_),
    .A2(_2265_),
    .B1(_2880_),
    .B2(_1672_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6899_ (.A1(_0975_),
    .A2(_2700_),
    .B1(_2881_),
    .B2(_2699_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6900_ (.A1(_2206_),
    .A2(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6901_ (.A1(_0976_),
    .A2(_2636_),
    .B1(_2878_),
    .B2(_2608_),
    .C(_2883_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6902_ (.A1(net50),
    .A2(_2794_),
    .B(_2826_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6903_ (.A1(_2607_),
    .A2(_2884_),
    .B(_2885_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6904_ (.A1(_1529_),
    .A2(_2861_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6905_ (.A1(_1529_),
    .A2(_2869_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6906_ (.A1(_2648_),
    .A2(_2886_),
    .B1(_2887_),
    .B2(_1827_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6907_ (.A1(net50),
    .A2(_2874_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6908_ (.A1(net37),
    .A2(_2889_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6909_ (.A1(_2693_),
    .A2(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6910_ (.A1(_2769_),
    .A2(_2888_),
    .B(_2891_),
    .C(_1821_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6911_ (.A1(_0975_),
    .A2(_1322_),
    .B(_2855_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6912_ (.A1(_2302_),
    .A2(_2893_),
    .B(_1788_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6913_ (.A1(_2302_),
    .A2(_2893_),
    .B(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6914_ (.A1(_1729_),
    .A2(_1818_),
    .A3(_2892_),
    .A4(_2895_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6915_ (.A1(_1760_),
    .A2(_2890_),
    .B(_2310_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6916_ (.A1(_1241_),
    .A2(_2665_),
    .B1(_2897_),
    .B2(_2790_),
    .C(_1939_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6917_ (.A1(_0980_),
    .A2(_2698_),
    .B1(_2898_),
    .B2(_2306_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6918_ (.A1(_2896_),
    .A2(_2899_),
    .B(_2705_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6919_ (.A1(net37),
    .A2(_2607_),
    .B(_1151_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6920_ (.A1(_2900_),
    .A2(_2901_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6921_ (.A1(net37),
    .A2(net50),
    .A3(_2874_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6922_ (.A1(net38),
    .A2(_2902_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6923_ (.A1(_2612_),
    .A2(_2903_),
    .B(_1847_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6924_ (.A1(_2858_),
    .A2(_2860_),
    .B(_1747_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6925_ (.A1(_2646_),
    .A2(_2390_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6926_ (.A1(_2866_),
    .A2(_2868_),
    .B(_1492_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6927_ (.I(_1494_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6928_ (.A1(_2908_),
    .A2(_2347_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6929_ (.A1(_2908_),
    .A2(_2905_),
    .B(_2907_),
    .C(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6930_ (.A1(_2905_),
    .A2(_2906_),
    .A3(_2907_),
    .B1(_2910_),
    .B2(_1535_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6931_ (.A1(_2814_),
    .A2(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6932_ (.A1(_2300_),
    .A2(_2301_),
    .A3(_2855_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6933_ (.A1(_2334_),
    .A2(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6934_ (.A1(_2333_),
    .A2(_2914_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6935_ (.A1(_2904_),
    .A2(_2912_),
    .B1(_2915_),
    .B2(_1857_),
    .C(_2457_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6936_ (.A1(_2667_),
    .A2(_2903_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6937_ (.A1(_1535_),
    .A2(_2139_),
    .B(_2917_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6938_ (.A1(_2666_),
    .A2(_2337_),
    .B1(_2918_),
    .B2(_2626_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6939_ (.A1(_1244_),
    .A2(_2665_),
    .B1(_2919_),
    .B2(_2623_),
    .C(_1582_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6940_ (.A1(_2916_),
    .A2(_2920_),
    .B(_1647_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6941_ (.A1(_1244_),
    .A2(_2637_),
    .B(_2921_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6942_ (.A1(net38),
    .A2(_2794_),
    .B(_2826_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6943_ (.A1(_2607_),
    .A2(_2922_),
    .B(_2923_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6944_ (.I(net38),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6945_ (.A1(_2924_),
    .A2(_2902_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6946_ (.A1(net39),
    .A2(_2925_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6947_ (.A1(_1494_),
    .A2(_2390_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6948_ (.A1(_2908_),
    .A2(_2905_),
    .B(_2907_),
    .C(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6949_ (.A1(_2389_),
    .A2(_2905_),
    .A3(_2906_),
    .A4(_2907_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6950_ (.A1(_1538_),
    .A2(_2928_),
    .B(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6951_ (.A1(_2814_),
    .A2(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6952_ (.A1(_1605_),
    .A2(_2926_),
    .B(_2931_),
    .C(_2638_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6953_ (.A1(_2333_),
    .A2(_2914_),
    .B(_2376_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6954_ (.A1(_2375_),
    .A2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6955_ (.A1(_1414_),
    .A2(_1296_),
    .B1(_2609_),
    .B2(_2934_),
    .C(_1755_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6956_ (.A1(_2211_),
    .A2(_2378_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6957_ (.A1(_1740_),
    .A2(_2926_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6958_ (.A1(_2382_),
    .A2(_2937_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6959_ (.A1(_1247_),
    .A2(_2787_),
    .B1(_2938_),
    .B2(_2790_),
    .C(_1887_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6960_ (.A1(_0989_),
    .A2(_2698_),
    .B1(_2932_),
    .B2(_2935_),
    .C1(_2936_),
    .C2(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6961_ (.A1(_2678_),
    .A2(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6962_ (.A1(net39),
    .A2(_2674_),
    .B(_1151_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6963_ (.A1(_2941_),
    .A2(_2942_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6964_ (.A1(net39),
    .A2(_2925_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6965_ (.A1(net40),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6966_ (.A1(_1538_),
    .A2(_2646_),
    .B(_2928_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6967_ (.A1(_1542_),
    .A2(_2929_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6968_ (.A1(_1542_),
    .A2(_2945_),
    .B(_2946_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6969_ (.A1(_2908_),
    .A2(_2944_),
    .B(_2947_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6970_ (.A1(_2404_),
    .A2(_2913_),
    .B(_2406_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6971_ (.A1(_2408_),
    .A2(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6972_ (.A1(_2814_),
    .A2(_2944_),
    .B1(_2950_),
    .B2(_1821_),
    .C(_2479_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6973_ (.A1(_1600_),
    .A2(_2948_),
    .B(_2951_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6974_ (.A1(_1740_),
    .A2(_2944_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6975_ (.A1(_2420_),
    .A2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6976_ (.A1(_1249_),
    .A2(_2787_),
    .B1(_2954_),
    .B2(_1443_),
    .C(_2410_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6977_ (.A1(_0993_),
    .A2(_2636_),
    .B1(_2955_),
    .B2(_1939_),
    .C(_2606_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6978_ (.A1(_1690_),
    .A2(_2952_),
    .B(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6979_ (.A1(net40),
    .A2(_2674_),
    .B(_0885_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6980_ (.A1(_2957_),
    .A2(_2958_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6981_ (.I(_3238_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6982_ (.I(_2959_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6983_ (.I(_2959_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6984_ (.A1(_2961_),
    .A2(_2462_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6985_ (.A1(_3317_),
    .A2(_2960_),
    .B(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6986_ (.A1(_1820_),
    .A2(_1415_),
    .B(_1143_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6987_ (.A1(_3171_),
    .A2(_1015_),
    .A3(_1604_),
    .A4(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6988_ (.A1(_1613_),
    .A2(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6989_ (.A1(_1011_),
    .A2(_1584_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6990_ (.A1(_1561_),
    .A2(_2437_),
    .A3(_2966_),
    .A4(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6991_ (.I(_2968_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6992_ (.I(_2968_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6993_ (.A1(net41),
    .A2(_2970_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6994_ (.A1(_2963_),
    .A2(_2969_),
    .B(_2971_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6995_ (.I(_2959_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_3494_),
    .A2(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6997_ (.A1(_2960_),
    .A2(_1118_),
    .B(_2973_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6998_ (.A1(net42),
    .A2(_2970_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6999_ (.A1(_2969_),
    .A2(_2974_),
    .B(_2975_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7000_ (.I(_2959_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7001_ (.A1(_2972_),
    .A2(_0726_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7002_ (.A1(_1713_),
    .A2(_2976_),
    .B(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7003_ (.A1(net43),
    .A2(_2970_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7004_ (.A1(_2969_),
    .A2(_2978_),
    .B(_2979_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7005_ (.A1(_2972_),
    .A2(_0741_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7006_ (.A1(_0725_),
    .A2(_2976_),
    .B(_2980_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7007_ (.A1(net44),
    .A2(_2970_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7008_ (.A1(_2969_),
    .A2(_2981_),
    .B(_2982_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7009_ (.I(_2968_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7010_ (.A1(_2972_),
    .A2(_0472_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7011_ (.A1(_0363_),
    .A2(_2976_),
    .B(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7012_ (.I(_2968_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7013_ (.A1(net45),
    .A2(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7014_ (.A1(_2983_),
    .A2(_2985_),
    .B(_2987_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7015_ (.A1(_2961_),
    .A2(_0772_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7016_ (.A1(_0471_),
    .A2(_2976_),
    .B(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7017_ (.A1(net19),
    .A2(_2986_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7018_ (.A1(_2983_),
    .A2(_2989_),
    .B(_2990_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7019_ (.A1(_2961_),
    .A2(_0785_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7020_ (.A1(_1728_),
    .A2(_2960_),
    .B(_2991_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7021_ (.A1(net20),
    .A2(_2986_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7022_ (.A1(_2983_),
    .A2(_2992_),
    .B(_2993_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7023_ (.A1(_2961_),
    .A2(_1141_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7024_ (.A1(_0585_),
    .A2(_2960_),
    .B(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7025_ (.A1(net21),
    .A2(_2986_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7026_ (.A1(_2983_),
    .A2(_2995_),
    .B(_2996_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7027_ (.A1(_3285_),
    .A2(_0798_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7028_ (.I(_2997_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7029_ (.A1(_3284_),
    .A2(_0798_),
    .B(_3449_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7030_ (.I(_2999_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7031_ (.A1(\as2650.r123[0][0] ),
    .A2(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7032_ (.A1(_3448_),
    .A2(_2998_),
    .B(_3001_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7033_ (.A1(\as2650.r123[0][1] ),
    .A2(_3000_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7034_ (.A1(_3530_),
    .A2(_2998_),
    .B(_3002_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7035_ (.A1(\as2650.r123[0][2] ),
    .A2(_3000_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7036_ (.A1(_0279_),
    .A2(_2998_),
    .B(_3003_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7037_ (.A1(\as2650.r123[0][3] ),
    .A2(_3000_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7038_ (.A1(_0354_),
    .A2(_2998_),
    .B(_3004_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7039_ (.I(_2997_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7040_ (.I(_2999_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7041_ (.A1(\as2650.r123[0][4] ),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7042_ (.A1(_0424_),
    .A2(_3005_),
    .B(_3007_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7043_ (.A1(\as2650.r123[0][5] ),
    .A2(_3006_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7044_ (.A1(_0499_),
    .A2(_3005_),
    .B(_3008_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7045_ (.A1(\as2650.r123[0][6] ),
    .A2(_3006_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7046_ (.A1(_0554_),
    .A2(_3005_),
    .B(_3009_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7047_ (.A1(\as2650.r123[0][7] ),
    .A2(_3006_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7048_ (.A1(_0605_),
    .A2(_3005_),
    .B(_3010_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7049_ (.A1(_3171_),
    .A2(_1307_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7050_ (.A1(_1573_),
    .A2(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7051_ (.A1(_1537_),
    .A2(_3011_),
    .B(_3012_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7052_ (.A1(_1567_),
    .A2(_3011_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7053_ (.A1(_1541_),
    .A2(_3011_),
    .B(_3013_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7054_ (.A1(_1566_),
    .A2(_0854_),
    .A3(_1653_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7055_ (.A1(_0671_),
    .A2(_1107_),
    .A3(_0827_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7056_ (.A1(_3479_),
    .A2(_1026_),
    .B(_1559_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7057_ (.A1(_1036_),
    .A2(_1019_),
    .A3(_3015_),
    .A4(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7058_ (.A1(_3229_),
    .A2(_0802_),
    .A3(_1055_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7059_ (.A1(_1009_),
    .A2(_3017_),
    .A3(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7060_ (.A1(_1060_),
    .A2(_3019_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7061_ (.A1(_1833_),
    .A2(_1578_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7062_ (.A1(_0853_),
    .A2(_1099_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7063_ (.A1(_3350_),
    .A2(_0637_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7064_ (.A1(_3326_),
    .A2(_3023_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7065_ (.A1(_1428_),
    .A2(_1041_),
    .B(_1015_),
    .C(_1145_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7066_ (.A1(_3022_),
    .A2(_3024_),
    .A3(_3025_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7067_ (.A1(_1012_),
    .A2(_3020_),
    .A3(_3021_),
    .A4(_3026_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7068_ (.A1(_0873_),
    .A2(_3014_),
    .B(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7069_ (.I(_0870_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7070_ (.A1(_0804_),
    .A2(_3029_),
    .B(_1726_),
    .C(_0808_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7071_ (.A1(_2539_),
    .A2(_2540_),
    .A3(_3030_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7072_ (.A1(_1094_),
    .A2(_0423_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7073_ (.A1(_1567_),
    .A2(_3031_),
    .B(_3028_),
    .C(_3032_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7074_ (.A1(_1178_),
    .A2(_3028_),
    .B(_3033_),
    .C(_2736_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7075_ (.A1(_1305_),
    .A2(_3014_),
    .B(_3027_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7076_ (.A1(_1700_),
    .A2(_0785_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7077_ (.A1(_0501_),
    .A2(_1701_),
    .B(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7078_ (.A1(_1700_),
    .A2(_0567_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7079_ (.A1(_0560_),
    .A2(_1701_),
    .B(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7080_ (.A1(_1700_),
    .A2(_0374_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7081_ (.A1(_0440_),
    .A2(_1701_),
    .B(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7082_ (.A1(_0299_),
    .A2(_0306_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7083_ (.A1(_3455_),
    .A2(_3483_),
    .B(_3439_),
    .C(_3445_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7084_ (.A1(_3580_),
    .A2(_1022_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7085_ (.A1(_1022_),
    .A2(_3504_),
    .B(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7086_ (.A1(_3455_),
    .A2(_1086_),
    .B1(_0277_),
    .B2(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7087_ (.A1(_0277_),
    .A2(_3044_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7088_ (.A1(_0299_),
    .A2(_0306_),
    .B1(_3042_),
    .B2(_3045_),
    .C(_3046_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7089_ (.A1(_0418_),
    .A2(_0422_),
    .B1(_3041_),
    .B2(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7090_ (.A1(_0418_),
    .A2(_0422_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7091_ (.A1(_0452_),
    .A2(_3040_),
    .B(_3048_),
    .C(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7092_ (.A1(_0453_),
    .A2(_3040_),
    .B1(_0527_),
    .B2(_3036_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7093_ (.A1(_3050_),
    .A2(_3051_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7094_ (.A1(_0528_),
    .A2(_3036_),
    .B1(_1085_),
    .B2(_3038_),
    .C(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7095_ (.A1(_0577_),
    .A2(_3038_),
    .B(_1204_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7096_ (.A1(_1128_),
    .A2(_2018_),
    .A3(_0804_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7097_ (.A1(_1698_),
    .A2(_3055_),
    .B(_2465_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7098_ (.A1(_2465_),
    .A2(_0773_),
    .B(_3056_),
    .C(_2471_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7099_ (.A1(_2471_),
    .A2(_2462_),
    .B(_3057_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7100_ (.A1(_3053_),
    .A2(_3054_),
    .B1(_3058_),
    .B2(_1759_),
    .C(_3034_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7101_ (.A1(_3346_),
    .A2(_3034_),
    .B(_3059_),
    .C(_2736_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7102_ (.A1(_1085_),
    .A2(_3038_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7103_ (.A1(_1582_),
    .A2(_0559_),
    .A3(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7104_ (.A1(_0637_),
    .A2(_1555_),
    .A3(_3022_),
    .A4(_3025_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7105_ (.A1(_3193_),
    .A2(_1715_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7106_ (.A1(_1755_),
    .A2(_3063_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7107_ (.A1(_3020_),
    .A2(_3062_),
    .A3(_3064_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7108_ (.A1(_1713_),
    .A2(_1696_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7109_ (.A1(_0823_),
    .A2(_0805_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7110_ (.A1(_3066_),
    .A2(_3067_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7111_ (.A1(_1759_),
    .A2(_1715_),
    .A3(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7112_ (.A1(_3065_),
    .A2(_3069_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7113_ (.A1(\as2650.overflow ),
    .A2(_3065_),
    .B(_0884_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7114_ (.A1(_3061_),
    .A2(_3070_),
    .B(_3071_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7115_ (.I(_1125_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7116_ (.A1(_1570_),
    .A2(_1761_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7117_ (.A1(_1675_),
    .A2(_0878_),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7118_ (.A1(_1002_),
    .A2(_0831_),
    .A3(_1056_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7119_ (.A1(_1642_),
    .A2(_0829_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7120_ (.A1(_3073_),
    .A2(_3074_),
    .A3(_3075_),
    .A4(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7121_ (.A1(_3072_),
    .A2(_1697_),
    .B(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7122_ (.A1(_3072_),
    .A2(_0875_),
    .A3(_0805_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7123_ (.A1(_3073_),
    .A2(_3074_),
    .A3(_3075_),
    .A4(_3076_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7124_ (.A1(_1723_),
    .A2(_3079_),
    .B(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7125_ (.A1(_3258_),
    .A2(_3078_),
    .B(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7126_ (.A1(_2249_),
    .A2(_3082_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7127_ (.I(_1735_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7128_ (.I(_1132_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_1696_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7130_ (.A1(_3084_),
    .A2(_3085_),
    .B(_3077_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7131_ (.A1(_3084_),
    .A2(_0823_),
    .A3(_0805_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7132_ (.A1(_1720_),
    .A2(_3087_),
    .B(_3080_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7133_ (.A1(_3326_),
    .A2(_3086_),
    .B(_3088_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7134_ (.A1(_3083_),
    .A2(_3089_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7135_ (.A1(_1313_),
    .A2(_3085_),
    .B(_3077_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7136_ (.A1(_1064_),
    .A2(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7137_ (.A1(_0798_),
    .A2(_0878_),
    .A3(_1709_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7138_ (.A1(_1710_),
    .A2(_3077_),
    .A3(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7139_ (.A1(_3091_),
    .A2(_3093_),
    .B(_1794_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7140_ (.A1(_1165_),
    .A2(_0877_),
    .B(_1810_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7141_ (.A1(_0840_),
    .A2(_1861_),
    .A3(_0843_),
    .A4(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7143_ (.A1(_1322_),
    .A2(_0876_),
    .A3(_1729_),
    .A4(_0878_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7144_ (.A1(_1728_),
    .A2(_1714_),
    .B(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7145_ (.A1(_1546_),
    .A2(_1729_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(_3095_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7147_ (.A1(_3099_),
    .A2(_3100_),
    .B(net27),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7148_ (.A1(_3096_),
    .A2(_3098_),
    .B(_3101_),
    .C(_2736_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7149_ (.I(_3095_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7150_ (.A1(_3072_),
    .A2(_3085_),
    .B(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7151_ (.A1(_0876_),
    .A2(_0877_),
    .B(_1707_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_3104_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7153_ (.A1(_3072_),
    .A2(_3105_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7154_ (.A1(_1723_),
    .A2(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7155_ (.A1(\as2650.psu[4] ),
    .A2(_3103_),
    .B1(_3107_),
    .B2(_3096_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7156_ (.A1(_3083_),
    .A2(_3108_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7157_ (.A1(_3084_),
    .A2(_3085_),
    .B(_3102_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7158_ (.A1(_3084_),
    .A2(_3105_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7159_ (.A1(_1720_),
    .A2(_3110_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7160_ (.A1(\as2650.psu[3] ),
    .A2(_3109_),
    .B1(_3111_),
    .B2(_3096_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7161_ (.A1(_3083_),
    .A2(_3112_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7162_ (.A1(_1715_),
    .A2(_3100_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7163_ (.A1(_1130_),
    .A2(_3105_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7164_ (.A1(_3066_),
    .A2(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7165_ (.A1(\as2650.psu[2] ),
    .A2(_3113_),
    .B1(_3115_),
    .B2(_3096_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7166_ (.A1(_3083_),
    .A2(_3116_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7167_ (.A1(_1313_),
    .A2(_1643_),
    .B(_3102_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7168_ (.A1(_1313_),
    .A2(_3105_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7169_ (.A1(_1709_),
    .A2(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7170_ (.A1(\as2650.psu[1] ),
    .A2(_3117_),
    .B1(_3119_),
    .B2(_3100_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7171_ (.A1(_1794_),
    .A2(_3120_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7172_ (.A1(_1305_),
    .A2(_1643_),
    .B(_3102_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7173_ (.A1(_1305_),
    .A2(_3104_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7174_ (.A1(_1698_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7175_ (.A1(\as2650.psu[0] ),
    .A2(_3121_),
    .B1(_3123_),
    .B2(_3100_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7176_ (.A1(_1794_),
    .A2(_3124_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7177_ (.D(_0000_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7178_ (.D(_0001_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7179_ (.D(_0002_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7180_ (.D(_0003_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7181_ (.D(_0004_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7182_ (.D(_0005_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7183_ (.D(_0006_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7184_ (.D(_0007_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7185_ (.D(_0008_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7186_ (.D(_0009_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7187_ (.D(_0010_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7188_ (.D(_0011_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7189_ (.D(_0012_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7190_ (.D(_0013_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7191_ (.D(_0014_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7192_ (.D(_0015_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7193_ (.D(_0016_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7194_ (.D(_0017_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7195_ (.D(_0018_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7196_ (.D(_0019_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7197_ (.D(_0020_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7198_ (.D(_0021_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7199_ (.D(_0022_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7200_ (.D(_0023_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7201_ (.D(_0024_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7202_ (.D(_0025_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7203_ (.D(_0026_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7204_ (.D(_0027_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7205_ (.D(_0028_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7206_ (.D(_0029_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7207_ (.D(_0030_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7208_ (.D(_0031_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7209_ (.D(_0032_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7210_ (.D(_0033_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7211_ (.D(_0034_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7212_ (.D(_0035_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7213_ (.D(_0036_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7214_ (.D(_0037_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7215_ (.D(_0038_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7216_ (.D(_0039_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7217_ (.D(_0040_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7218_ (.D(_0041_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7219_ (.D(_0042_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7220_ (.D(_0043_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7221_ (.D(_0044_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7222_ (.D(_0045_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7223_ (.D(_0046_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7224_ (.D(_0047_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7225_ (.D(_0048_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7226_ (.D(_0049_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7227_ (.D(_0050_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7228_ (.D(_0051_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7229_ (.D(_0052_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7230_ (.D(_0053_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7231_ (.D(_0054_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7232_ (.D(_0055_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7233_ (.D(_0056_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7234_ (.D(_0057_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7235_ (.D(_0058_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7236_ (.D(_0059_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7237_ (.D(_0060_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7238_ (.D(_0061_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7239_ (.D(_0062_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7240_ (.D(_0063_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7241_ (.D(_0064_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7242_ (.D(_0065_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7243_ (.D(_0066_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7244_ (.D(_0067_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7245_ (.D(_0068_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7246_ (.D(_0069_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7247_ (.D(_0070_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7248_ (.D(_0071_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7249_ (.D(_0072_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7250_ (.D(_0073_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7251_ (.D(_0074_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7252_ (.D(_0075_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7253_ (.D(_0076_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7254_ (.D(_0077_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7255_ (.D(_0078_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7256_ (.D(_0079_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7257_ (.D(_0080_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7258_ (.D(_0081_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7259_ (.D(_0082_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7260_ (.D(_0083_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7261_ (.D(_0084_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7262_ (.D(_0085_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7263_ (.D(_0086_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7264_ (.D(_0087_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7265_ (.D(_0088_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7266_ (.D(_0089_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7267_ (.D(_0090_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7268_ (.D(_0091_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7269_ (.D(_0092_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7270_ (.D(_0093_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7271_ (.D(_0094_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7272_ (.D(_0095_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7273_ (.D(_0096_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7274_ (.D(_0097_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7275_ (.D(_0098_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7276_ (.D(_0099_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7277_ (.D(_0100_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7278_ (.D(_0101_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7279_ (.D(_0102_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7280_ (.D(_0103_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7281_ (.D(_0104_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7282_ (.D(_0105_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7283_ (.D(_0106_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7284_ (.D(_0107_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7285_ (.D(_0108_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7286_ (.D(_0109_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7287_ (.D(_0110_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7288_ (.D(_0111_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7289_ (.D(_0112_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7290_ (.D(_0113_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7291_ (.D(_0114_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7292_ (.D(_0115_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7293_ (.D(_0116_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7294_ (.D(_0117_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7295_ (.D(_0118_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7296_ (.D(_0119_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7297_ (.D(_0120_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7298_ (.D(_0121_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7299_ (.D(_0122_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7300_ (.D(_0123_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7301_ (.D(_0124_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7302_ (.D(_0125_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7303_ (.D(_0126_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7304_ (.D(_0127_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7305_ (.D(_0128_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7306_ (.D(_0129_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7307_ (.D(_0130_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7308_ (.D(_0131_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7309_ (.D(_0132_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7310_ (.D(_0133_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7311_ (.D(_0134_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7312_ (.D(_0135_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7313_ (.D(_0136_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7314_ (.D(_0137_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7315_ (.D(_0138_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7316_ (.D(_0139_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7317_ (.D(_0140_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7318_ (.D(_0141_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7319_ (.D(_0142_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7320_ (.D(_0143_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7321_ (.D(_0144_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7322_ (.D(_0145_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7323_ (.D(_0146_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7324_ (.D(_0147_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7325_ (.D(_0148_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7326_ (.D(_0149_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7327_ (.D(_0150_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7328_ (.D(_0151_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7329_ (.D(_0152_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7330_ (.D(_0153_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7331_ (.D(_0154_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7332_ (.D(_0155_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7333_ (.D(_0156_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7334_ (.D(_0157_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7335_ (.D(_0158_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7336_ (.D(_0159_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7337_ (.D(_0160_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7338_ (.D(_0161_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7339_ (.D(_0162_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7340_ (.D(_0163_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7341_ (.D(_0164_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7342_ (.D(_0165_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7343_ (.D(_0166_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7344_ (.D(_0167_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7345_ (.D(_0168_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7346_ (.D(_0169_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7347_ (.D(_0170_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7348_ (.D(_0171_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7349_ (.D(_0172_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7350_ (.D(_0173_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7351_ (.D(_0174_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7352_ (.D(_0175_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7353_ (.D(_0176_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7354_ (.D(_0177_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7355_ (.D(_0178_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7356_ (.D(_0179_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7357_ (.D(_0180_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7358_ (.D(_0181_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7359_ (.D(_0182_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7360_ (.D(_0183_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7361_ (.D(_0184_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7362_ (.D(_0185_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7363_ (.D(_0186_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7364_ (.D(_0187_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7365_ (.D(_0188_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7366_ (.D(_0189_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7367_ (.D(_0190_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7368_ (.D(_0191_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7369_ (.D(_0192_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7370_ (.D(_0193_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7371_ (.D(_0194_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7372_ (.D(_0195_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7373_ (.D(_0196_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7374_ (.D(_0197_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7375_ (.D(_0198_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7376_ (.D(_0199_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7377_ (.D(_0200_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7378_ (.D(_0201_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7379_ (.D(_0202_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7380_ (.D(_0203_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7381_ (.D(_0204_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7382_ (.D(_0205_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7383_ (.D(_0206_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7384_ (.D(_0207_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7385_ (.D(_0208_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7386_ (.D(_0209_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7387_ (.D(_0210_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7388_ (.D(_0211_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7389_ (.D(_0212_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7390_ (.D(_0213_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7391_ (.D(_0214_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7392_ (.D(_0215_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7393_ (.D(_0216_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7394_ (.D(_0217_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7395_ (.D(_0218_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7396_ (.D(_0219_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7397_ (.D(_0220_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7398_ (.D(_0221_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7399_ (.D(_0222_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7400_ (.D(_0223_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7401_ (.D(_0224_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7402_ (.D(_0225_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7403_ (.D(_0226_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7404_ (.D(_0227_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7405_ (.D(_0228_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7406_ (.D(_0229_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7407_ (.D(_0230_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7408_ (.D(_0231_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7409_ (.D(_0232_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7410_ (.D(_0233_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7411_ (.D(_0234_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7412_ (.D(_0235_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7413_ (.D(_0236_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7414_ (.D(_0237_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7415_ (.D(_0238_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7416_ (.D(_0239_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7417_ (.D(_0240_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7418_ (.D(_0241_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7419_ (.D(_0242_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7420_ (.D(_0243_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7421_ (.D(_0244_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7422_ (.D(_0245_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7423_ (.D(_0246_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7424_ (.D(_0247_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7425_ (.D(_0248_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7426_ (.D(_0249_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7427_ (.D(_0250_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7428_ (.D(_0251_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7429_ (.D(_0252_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7430_ (.D(_0253_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7431_ (.D(_0254_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7432_ (.D(_0255_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7433_ (.D(_0256_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7434_ (.D(_0257_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7435_ (.D(_0258_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7436_ (.D(_0259_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7437_ (.D(_0260_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7479_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7480_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7481_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7482_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7483_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7484_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7485_ (.I(net47),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(io_in[5]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[6]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[7]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net49),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net52),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net51),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net13),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net36),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net33),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net29),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout53 (.I(net26),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__D (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__D (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__D (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__D (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__D (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__D (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__D (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__D (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__D (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__B1 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__I (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A3 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__B (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__B2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__B1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__I (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A3 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I0 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__I1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A4 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__B (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__B (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__B (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__I (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__B2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__C (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__B (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__B (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A4 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__I (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__B (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A3 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__I (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__C1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A3 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__B2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__I (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__B (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__I (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__C1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__B (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__C2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__B2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__B2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__B2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A3 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__B (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__C (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__B1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__C (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__I1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__I (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A3 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__I (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__B (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__I1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__B1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__B (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A4 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A3 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A3 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__B1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A4 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__C (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A3 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A3 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__B2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I0 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__I (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__C1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__C2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__B (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__S (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__B (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__I (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A3 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__B1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A2 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__I (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__B (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__B1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__C1 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__B (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__B2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A3 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__B (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A4 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__C (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__I (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__B (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__I (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A3 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__B (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A4 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A3 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A3 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A3 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A4 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A3 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__C (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I0 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__I0 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I0 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A3 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__S (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__S (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__B (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__B1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A3 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__B (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A4 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__B (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__B1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__I1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A2 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I0 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I0 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I0 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A3 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A3 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A3 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__C (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__B (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__C (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__B (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__B (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__I (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A3 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__I (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__I (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__I (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__C (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A4 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__C (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__B (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__C (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A3 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__S (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A3 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__B (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A3 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__I (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__I (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__B (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A3 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__C (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A3 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__B (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A4 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__B (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A3 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__B (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A3 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A4 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A3 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__B (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__B (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__B (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__B (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__B (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__B2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__B2 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__B2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__S1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__B (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__B2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__B (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__I (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__B (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__B1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A4 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A3 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A4 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A4 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A3 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__I (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A3 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__S0 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__S0 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__B2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__B2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__B (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A3 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__I (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__S (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__I (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__I (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__I (.I(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__I0 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__I0 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I0 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__I0 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A3 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__I (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A2 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A3 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A3 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A3 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__B2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__B (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__B1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A3 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__C (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A3 (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__B2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__C (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__B (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__B (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__B (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A3 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__B1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__B (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A3 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A3 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A4 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A3 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A4 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A4 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__B (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__I (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__B (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__B (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A3 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A2 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A3 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__C (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__I (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__C (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A3 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A3 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A3 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__S (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__B (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A3 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__B (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__I (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__B2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__C (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__B (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__B (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__I (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__B (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__C (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__B (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__I (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__B2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__C (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__C (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__C (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__C (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__C (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__B (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A3 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__B (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__I (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__C (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__C (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__C (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A3 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__B2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A3 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A4 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__B (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__C (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__C (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__B1 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__B (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A3 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__C (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__I (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__B (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__C (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__B (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__B (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__C (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__C (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__I (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__C (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__C (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__B (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__C (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__B2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A3 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A3 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__C (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__I (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__B1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__B1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__B2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A2 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__B1 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A4 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A3 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__C (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__B (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__B1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__B2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__B2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A3 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__S (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__S (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__S (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__S (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__S (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__I1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__C (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A2 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__I1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__S (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__S (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__S (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__S (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__I1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__I1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I0 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I0 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__I1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__S (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__S (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__S (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__S (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__I1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__I1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__I1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__S (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__S (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__S (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__S (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__S (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__S (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__S (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__S (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__S (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__S (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__S (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__S (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__S (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__S (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__I (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A3 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__B (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__I (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A4 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__C (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__B1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__B1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__B1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__B2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__C (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__B2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I0 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__B2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__S (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__S (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__I (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__I (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__S (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__S (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__S (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__B2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__C (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__B (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A3 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__B (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A3 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__B2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__B (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__B2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__C (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__C (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A3 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__I (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__I (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__B (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__B (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__B (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__B2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A4 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__C (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__C (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__B2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__C (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A1 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__I (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__I (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__C (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__B2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__C (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__C (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__C (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__C (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__I (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__C (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__S (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__S (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A4 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__B (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__C (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A3 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A3 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__B1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__B2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A3 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__C (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__C (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__B (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__B (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__B1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__C (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__S (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__B2 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__I (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__B2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__I (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__I (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A3 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__B1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__B (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__I (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__B1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__B (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__B2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__C (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__B2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__B (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__I (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__C (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__C (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__C (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__C (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__C (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__B (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A4 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__B (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__C (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__C (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A3 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A4 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__C (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__C (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__C (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__B (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__C (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__B (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__B (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__C (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__B2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__B1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A3 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A3 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A4 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A4 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A3 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__C (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A4 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A4 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__B2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__C (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__B (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__B (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A4 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A3 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A3 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__I (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__B (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__B (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__B (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__B (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__I (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__B2 (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__B (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__B (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__C (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__B (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A3 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__C (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__C (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__B (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A3 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__B1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__B1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A4 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A4 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A3 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__B (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__C (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__B (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__B2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__B2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A4 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A3 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__B (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A3 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__B (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__C (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__B2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__C (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__C (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__C (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__C (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__B (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__I0 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__S (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__S (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__S (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__S (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__S (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__S (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__B (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__B2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__B (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A3 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__B (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I0 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__B (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__B2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__I (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A3 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__B (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I0 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__B (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I0 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__B (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__I0 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A3 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__I0 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__B (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__I (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__C (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__C (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__B (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__B (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__B (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A4 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__C (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__C (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__C (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__C (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__C (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__C (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__B2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__B2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__B (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I (.I(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__B (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A2 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__C (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A3 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__B2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__B (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__B2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__C (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__C (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__B (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__B2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A3 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__C (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__B (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__B (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__B (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__B (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__C (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__C (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__B (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__B2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__I (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__B2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__B (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A3 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__B2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__B (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__C (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__B1 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A4 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__B2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__C (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__B2 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__C (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A3 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__B (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A2 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__C (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__C (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__C (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__B2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__B (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__B1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__B2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__B (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__B (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__C2 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A3 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A4 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__B2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__I (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__B2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__B2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A1 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A3 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A3 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A4 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A3 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A3 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__C (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__I (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__I (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__C (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__I (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__B2 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__I (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A3 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__I (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__B1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__I (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__I (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__B1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__B (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__C (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__B2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__B1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__B2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__B1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__B1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__B1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__B2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__B2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__C (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__B2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__B2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__B2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__B2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__B2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A2 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__B2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__C (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__C (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__B1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__B1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__C (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__B (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__B (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__B1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__B2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__S0 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__B2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__B1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__I (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__B2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__B (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__C (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__C (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__C (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__C (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A3 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__B1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__B2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__B2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__B2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__B2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__B (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__B2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__B (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__C (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__C (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__C (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__B (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__B2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__B (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__B2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__B2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__B2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__B2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__B2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__B1 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__C (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__B (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__B (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__C (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__C (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__C (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__C (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__B (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__B2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__B2 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__C (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__B (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__I (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__B (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__B1 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__B (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__B1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__C (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__B (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__S1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__B2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__C (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__B1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__B2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__C (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__C (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__C (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__C (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__C (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__B1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__B1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__C (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__B (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__B2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__B1 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__B2 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__B2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__B2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__B2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__B2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__C (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__B (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A3 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__B (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A3 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__B2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__B2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__B2 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__S1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__B1 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__B2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__B2 (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__B (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__B1 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__C (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__B2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__B (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__C (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__C (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A3 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__B2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__I (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__B (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__B (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__B1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__B (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__B1 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__B2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__B (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A3 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__B2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__B (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__B (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__B1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__B1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__B2 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__B (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__B (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__B (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__B (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__B (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__B (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__B (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__B (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I0 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A3 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__B1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__B2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__I (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A3 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__B1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A3 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__B (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A3 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A4 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A3 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A3 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__C (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__C (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__B (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__B (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__C (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__I (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__C (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__C (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__C (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A3 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__C (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__C (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__B (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__B (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__B1 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__B (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__C (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A4 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__B (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__C (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A3 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__C (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__B (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__B (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__C (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A3 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__I (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__I (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__I (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__I (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__S (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__I (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__C (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__C (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__I (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__B2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__B2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__B2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A1 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__B1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__B (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__I (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A1 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A2 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__B (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__C (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__B (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__B (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__B1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__B2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__B2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__B2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__I (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__B2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__B2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__B2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__B2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__B1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__A2 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__I (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__I (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__C (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__B (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__I (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__B (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__C (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A2 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__I (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__B (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__B1 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__B (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__B2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A1 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A1 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A2 (.I(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A1 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A2 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__B (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A2 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__B1 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__B2 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__B2 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__B2 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__B2 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__B2 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__B (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__B (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__C (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__B2 (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A2 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A2 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A3 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A3 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__B (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__B (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__B1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__C (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__C (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__C (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__C (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A2 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A2 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A2 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A4 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A3 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A2 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__C (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__B (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__B (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__B (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__B (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A3 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A3 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A2 (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__A2 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A2 (.I(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__B (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A2 (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__B1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A2 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__B (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A2 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__B1 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A1 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__B (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A3 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__B (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A1 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A2 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__C (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A2 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__B (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A4 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A1 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A4 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__B (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A3 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__B (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A2 (.I(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__B1 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__B1 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__B1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__B1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__B (.I(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__I (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__I (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A2 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A2 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__I (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A3 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A4 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A3 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__B (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__B (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__B (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__C (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A2 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A3 (.I(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A3 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A3 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A2 (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__B (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__B (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__B (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__B (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__B (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A3 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__I (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__I (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__I (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__B2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__B2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__B (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__B2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__B2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__B (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__B (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__B (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__B (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__A2 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A2 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__S0 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A2 (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__I (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__I (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__C (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__I (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__S (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__S (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__S1 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__I (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__S1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__S (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__I (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__I (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__S (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__S (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__I (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__S (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__S (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__S (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__S (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__I (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__S0 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__S0 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__S0 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__S0 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__S0 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__I (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A3 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__I (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__I (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__I (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A3 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__I (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__I (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__I (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__I (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A3 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A1 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__B2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A3 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A2 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__I (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__I (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3648__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A2 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A2 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__I (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__I (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A3 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__I (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A3 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__I (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__I (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__I (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__B (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__A1 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A2 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A1 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A3 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3679__A4 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A2 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__A2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A3 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A4 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A3 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__B (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A3 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A3 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A3 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A3 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A3 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__I (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__B2 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A3 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A3 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A3 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__I (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A4 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A4 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A3 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__B (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A2 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A3 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__I (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A3 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A3 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__I (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A3 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A4 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A3 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__I (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__I (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__I (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__C (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__I (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__C (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__C (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__C (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__I (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A1 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__I (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__I (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A3 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A4 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__B (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__I (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__B1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A3 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__C (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__I (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__I (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A4 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A1 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__I (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__I (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__S (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__S1 (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__S (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A3 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A1 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__I (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__C1 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__C2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__B2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__B2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__I (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__B (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A3 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A3 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__I (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A1 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__B2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__S (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__I (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__B2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__I (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__I (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A4 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__A4 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__I (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A2 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3809__I (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A2 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__B (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A1 (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__B (.I(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A2 (.I(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__C (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__B (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__I (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__I (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A2 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__I (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__I (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__B1 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__A1 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__A2 (.I(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A3 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__I (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__I (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__I (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A3 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__I (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__I (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__B (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__I (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__B2 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__B2 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3857__I (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A3 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A1 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A1 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__C (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__C (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__I (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__I (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__C (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__I (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A1 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__I1 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__A1 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__B (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__C (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A1 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A1 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A2 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__B (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__I (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__I (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A1 (.I(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A1 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__I (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__B (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A3 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A2 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__C (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__I (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__C1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__C (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__B (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A1 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A1 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I1 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__S (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__S (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__S (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__B (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__B (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__B (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__A2 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I1 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A1 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A3 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__B (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__I (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__I (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A1 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A1 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__I (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__C (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__C (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__I (.I(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A3 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A2 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A2 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__S (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__S1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__S1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__S1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A3 (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A3 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__B (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__A1 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__B (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A1 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__I (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__B2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__I (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__I (.I(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A1 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__B2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A3 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A3 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__C (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__B (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A3 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A3 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A3 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A3 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A2 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A2 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A3 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A4 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A3 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A3 (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__B (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__B (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A1 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A3 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A2 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__A4 (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A3 (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A3 (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A4 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__I (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A4 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A2 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A4 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__I (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__I (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__B1 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__I (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__C (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__B (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A1 (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__I (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A3 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__C (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__I (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__I (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A2 (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__I (.I(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__A2 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A2 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__I (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A3 (.I(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__B2 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__I (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__B (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__B2 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__B2 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3754__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A4 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A3 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__I0 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I1 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__I0 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I1 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I1 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I1 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__I3 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__I1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__I3 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__I1 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I3 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__I1 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I3 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__I1 (.I(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__B1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__B1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I0 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I0 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I0 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I3 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__I3 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__I3 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__I (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__B1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__B (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__B (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__B2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A3 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__B (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__CLK (.I(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__CLK (.I(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__CLK (.I(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__CLK (.I(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__CLK (.I(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__CLK (.I(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__CLK (.I(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__CLK (.I(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net89;
 assign io_oeb[13] = net94;
 assign io_oeb[14] = net54;
 assign io_oeb[15] = net55;
 assign io_oeb[16] = net56;
 assign io_oeb[17] = net57;
 assign io_oeb[18] = net58;
 assign io_oeb[19] = net59;
 assign io_oeb[1] = net90;
 assign io_oeb[20] = net60;
 assign io_oeb[21] = net61;
 assign io_oeb[22] = net62;
 assign io_oeb[23] = net63;
 assign io_oeb[24] = net64;
 assign io_oeb[25] = net65;
 assign io_oeb[26] = net66;
 assign io_oeb[27] = net67;
 assign io_oeb[28] = net68;
 assign io_oeb[29] = net69;
 assign io_oeb[2] = net91;
 assign io_oeb[30] = net70;
 assign io_oeb[31] = net71;
 assign io_oeb[32] = net72;
 assign io_oeb[33] = net73;
 assign io_oeb[34] = net74;
 assign io_oeb[35] = net75;
 assign io_oeb[36] = net76;
 assign io_oeb[37] = net77;
 assign io_oeb[3] = net92;
 assign io_oeb[4] = net93;
 assign io_out[0] = net78;
 assign io_out[13] = net83;
 assign io_out[1] = net79;
 assign io_out[2] = net80;
 assign io_out[33] = net84;
 assign io_out[34] = net85;
 assign io_out[35] = net86;
 assign io_out[36] = net87;
 assign io_out[37] = net88;
 assign io_out[3] = net81;
 assign io_out[4] = net82;
endmodule

