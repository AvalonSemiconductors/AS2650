// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack_ptr[0] ;
 wire \as2650.stack_ptr[1] ;
 wire \as2650.stack_ptr[2] ;
 wire net89;
 wire clknet_leaf_1_wb_clk_i;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net90;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net91;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net92;
 wire net93;
 wire net78;
 wire net83;
 wire net79;
 wire net80;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net81;
 wire net82;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_1_1_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3940_ (.I(net26),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3941_ (.I(\as2650.psl[4] ),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3942_ (.I(_3477_),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3943_ (.I(_3478_),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3944_ (.I(_3479_),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3945_ (.I(_3480_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3946_ (.I(_3481_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3947_ (.I(_3482_),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3948_ (.I(_3483_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(\as2650.cycle[1] ),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3950_ (.I(\as2650.cycle[0] ),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3951_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3952_ (.A1(\as2650.cycle[3] ),
    .A2(\as2650.cycle[2] ),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3953_ (.A1(_3485_),
    .A2(_3486_),
    .A3(_3487_),
    .A4(_3488_),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3954_ (.I(_3489_),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3955_ (.I(_3490_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(\as2650.ins_reg[1] ),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3957_ (.I(_3492_),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3958_ (.I(_3493_),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3959_ (.I(_3494_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3960_ (.I(_3495_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3961_ (.I(_3496_),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3962_ (.I(\as2650.ins_reg[4] ),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3963_ (.I(_3498_),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3964_ (.I(\as2650.ins_reg[5] ),
    .Z(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3965_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3966_ (.I(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3967_ (.I(_3502_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3968_ (.A1(_3500_),
    .A2(_3503_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3969_ (.I(\as2650.ins_reg[6] ),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3970_ (.I(\as2650.ins_reg[7] ),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3971_ (.I(_3506_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3972_ (.A1(_3505_),
    .A2(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3973_ (.A1(_3499_),
    .A2(_3504_),
    .A3(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3974_ (.A1(_3497_),
    .A2(_3509_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(_3491_),
    .A2(_3510_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3976_ (.I(\as2650.halted ),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3977_ (.I(net10),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3978_ (.A1(_3512_),
    .A2(_3513_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3979_ (.I(_3514_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3980_ (.A1(_3484_),
    .A2(_3511_),
    .A3(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3981_ (.I(_3516_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3982_ (.I(_3517_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3983_ (.I(net10),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3984_ (.I(\as2650.ins_reg[0] ),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3985_ (.I(_3520_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3986_ (.I(_3521_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3987_ (.I(_3522_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3988_ (.A1(_3523_),
    .A2(_3495_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3989_ (.I(\as2650.cycle[1] ),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3990_ (.I(_3486_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3991_ (.I(_3487_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3992_ (.I(_3488_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3993_ (.A1(_3525_),
    .A2(_3526_),
    .A3(_3527_),
    .A4(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3994_ (.I(_3529_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3995_ (.I(\as2650.ins_reg[1] ),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3996_ (.I(_3531_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3997_ (.I(_3532_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3998_ (.I(_3533_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3999_ (.I(_3509_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4000_ (.A1(_3534_),
    .A2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4001_ (.A1(_3530_),
    .A2(_3536_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4002_ (.A1(_3482_),
    .A2(_3514_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4003_ (.A1(_3537_),
    .A2(_3538_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4004_ (.I(\as2650.ins_reg[4] ),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4005_ (.I(_3540_),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4006_ (.I(_3541_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4007_ (.I(_3542_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4008_ (.A1(_3485_),
    .A2(\as2650.cycle[0] ),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4009_ (.A1(_3527_),
    .A2(_3544_),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4010_ (.I(\as2650.cycle[2] ),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4011_ (.A1(\as2650.cycle[3] ),
    .A2(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4012_ (.A1(_3545_),
    .A2(_3547_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4013_ (.I(_3503_),
    .Z(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4014_ (.I(\as2650.ins_reg[0] ),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4015_ (.I(_3550_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4016_ (.A1(_3551_),
    .A2(_3533_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4017_ (.I(_3552_),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4018_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4019_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4020_ (.A1(_3554_),
    .A2(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4021_ (.I(\as2650.ins_reg[5] ),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4022_ (.I(\as2650.ins_reg[6] ),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4023_ (.I(\as2650.ins_reg[7] ),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4024_ (.A1(_3557_),
    .A2(_3558_),
    .A3(_3559_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4025_ (.A1(_3549_),
    .A2(_3553_),
    .A3(_3556_),
    .A4(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4026_ (.A1(_3543_),
    .A2(_3548_),
    .A3(_3561_),
    .ZN(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4027_ (.A1(_3538_),
    .A2(_3562_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4028_ (.A1(_3485_),
    .A2(\as2650.cycle[0] ),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4029_ (.A1(_3527_),
    .A2(_3528_),
    .A3(_3564_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4030_ (.I(\as2650.ins_reg[4] ),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4031_ (.A1(\as2650.ins_reg[3] ),
    .A2(_3566_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4032_ (.I(\as2650.ins_reg[2] ),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4033_ (.I(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4034_ (.A1(_3569_),
    .A2(_3557_),
    .A3(_3540_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4035_ (.A1(_3506_),
    .A2(_3570_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4036_ (.A1(_3565_),
    .A2(_3567_),
    .A3(_3571_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4037_ (.I(_3568_),
    .Z(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4038_ (.A1(_3558_),
    .A2(_3559_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4039_ (.A1(_3540_),
    .A2(_3574_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4040_ (.A1(_3573_),
    .A2(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4041_ (.A1(_3489_),
    .A2(_3567_),
    .A3(_3576_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4042_ (.I(_3507_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4043_ (.A1(\as2650.ins_reg[4] ),
    .A2(_3558_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4044_ (.A1(_3568_),
    .A2(_3500_),
    .A3(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4045_ (.I(_3580_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4046_ (.A1(_3578_),
    .A2(_3581_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4047_ (.A1(_3577_),
    .A2(_3582_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4048_ (.A1(_3572_),
    .A2(_3583_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4049_ (.I(_3499_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4050_ (.I(\as2650.cycle[7] ),
    .Z(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4051_ (.I(\as2650.cycle[5] ),
    .Z(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4052_ (.I(\as2650.cycle[4] ),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4053_ (.A1(_3485_),
    .A2(_3486_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4054_ (.A1(\as2650.cycle[6] ),
    .A2(_3528_),
    .A3(_3589_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4055_ (.A1(_3586_),
    .A2(_3587_),
    .A3(_3588_),
    .A4(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4056_ (.A1(_3585_),
    .A2(_3591_),
    .A3(_3556_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4057_ (.I(\as2650.ins_reg[3] ),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4058_ (.I(_3593_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4059_ (.I(_3559_),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4060_ (.A1(_3595_),
    .A2(_3580_),
    .ZN(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4061_ (.I(_3596_),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4062_ (.A1(_3594_),
    .A2(_3530_),
    .A3(_3597_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4063_ (.A1(_3592_),
    .A2(_3598_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4064_ (.I(\as2650.addr_buff[7] ),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4065_ (.A1(\as2650.cycle[5] ),
    .A2(_3588_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4066_ (.A1(\as2650.cycle[7] ),
    .A2(_3601_),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4067_ (.A1(_3590_),
    .A2(_3602_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4068_ (.A1(_3600_),
    .A2(_3603_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4069_ (.I(\as2650.addr_buff[6] ),
    .Z(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4070_ (.I(\as2650.addr_buff[5] ),
    .Z(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4071_ (.A1(_3605_),
    .A2(_3606_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4072_ (.A1(_3543_),
    .A2(_3607_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(_3604_),
    .A2(_3608_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4074_ (.A1(_3599_),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4075_ (.I(_3594_),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(_3611_),
    .A2(_3491_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4077_ (.A1(_3579_),
    .A2(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4078_ (.I(_3531_),
    .Z(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4079_ (.A1(_3520_),
    .A2(_3614_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4080_ (.I(_3615_),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4081_ (.I(_3616_),
    .Z(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4082_ (.I(_3617_),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4083_ (.A1(_3483_),
    .A2(_3514_),
    .A3(_3618_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4084_ (.I(_3619_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4085_ (.I(_3620_),
    .Z(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4086_ (.A1(_3584_),
    .A2(_3610_),
    .A3(_3613_),
    .B(_3621_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4087_ (.A1(_3568_),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4088_ (.I(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4089_ (.I(_3624_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4090_ (.A1(_3558_),
    .A2(_3559_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4091_ (.A1(_3500_),
    .A2(_3541_),
    .A3(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(_3625_),
    .A2(_3627_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4093_ (.A1(_3529_),
    .A2(_3628_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4094_ (.A1(_3620_),
    .A2(_3629_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4095_ (.I(_3630_),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4096_ (.I(_3631_),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4097_ (.A1(_3539_),
    .A2(_3563_),
    .A3(_3622_),
    .A4(_3632_),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4098_ (.A1(_3524_),
    .A2(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4099_ (.A1(_3519_),
    .A2(_3634_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4100_ (.I(_3635_),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4101_ (.I(_3631_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4102_ (.A1(_3538_),
    .A2(_3552_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4103_ (.A1(_3593_),
    .A2(_3596_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4104_ (.A1(_3489_),
    .A2(_3639_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4105_ (.A1(_3638_),
    .A2(_3640_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4106_ (.I(_3641_),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4107_ (.I(\as2650.psl[3] ),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4108_ (.I(_3643_),
    .Z(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4109_ (.I(\as2650.r0[7] ),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4110_ (.A1(_3480_),
    .A2(\as2650.r123_2[0][7] ),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4111_ (.I(_3477_),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4112_ (.I(_3647_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4113_ (.I(_3648_),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4114_ (.I(_3649_),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4115_ (.A1(_3650_),
    .A2(\as2650.r123[0][7] ),
    .B(_3495_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4116_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_3479_),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4117_ (.A1(_3533_),
    .A2(_3652_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4118_ (.A1(_3646_),
    .A2(_3651_),
    .B(_3653_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4119_ (.A1(_3480_),
    .A2(\as2650.r123[1][7] ),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4120_ (.A1(_3650_),
    .A2(\as2650.r123_2[1][7] ),
    .B(_3495_),
    .C(_3551_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4121_ (.A1(_3655_),
    .A2(_3656_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4122_ (.A1(_3645_),
    .A2(_3617_),
    .B1(_3654_),
    .B2(_3523_),
    .C(_3657_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4123_ (.I(_3658_),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4124_ (.I(_3659_),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4125_ (.I(_3660_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4126_ (.A1(_3643_),
    .A2(\as2650.carry ),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4127_ (.I(_3662_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4128_ (.A1(_3644_),
    .A2(_3661_),
    .B(_3663_),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4129_ (.I(net5),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4130_ (.I(_3665_),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4131_ (.I(_3666_),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4132_ (.A1(_3638_),
    .A2(_3572_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4133_ (.I(_3668_),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4134_ (.A1(_3667_),
    .A2(_3669_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4135_ (.I(_3487_),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4136_ (.I(_3488_),
    .Z(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4137_ (.A1(_3671_),
    .A2(_3672_),
    .A3(_3564_),
    .ZN(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4138_ (.I(_3567_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4139_ (.I(_3571_),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4140_ (.A1(_3674_),
    .A2(_3675_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4141_ (.A1(_3673_),
    .A2(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(_3620_),
    .A2(_3677_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4143_ (.A1(_3498_),
    .A2(_3505_),
    .A3(_3506_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4144_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123_2[1][0] ),
    .S(\as2650.psl[4] ),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4145_ (.I(\as2650.r0[0] ),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4146_ (.A1(_3681_),
    .A2(_3531_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4147_ (.A1(_3532_),
    .A2(_3680_),
    .B(_3682_),
    .C(_3550_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4148_ (.I(\as2650.r123_2[0][0] ),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4149_ (.I0(\as2650.r123[0][0] ),
    .I1(_3684_),
    .I2(\as2650.r123[2][0] ),
    .I3(\as2650.r123_2[2][0] ),
    .S0(\as2650.psl[4] ),
    .S1(_3531_),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(\as2650.ins_reg[0] ),
    .A2(_3685_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4151_ (.A1(_3683_),
    .A2(_3686_),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4152_ (.I(_3687_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4153_ (.I(_3688_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4154_ (.I(_3689_),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4155_ (.I(_3690_),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4156_ (.A1(_3679_),
    .A2(_3691_),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4157_ (.I(_3638_),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4158_ (.A1(_3693_),
    .A2(_3583_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4159_ (.I(_3694_),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4160_ (.A1(_3678_),
    .A2(_3692_),
    .B(_3695_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4161_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123_2[1][1] ),
    .S(_3477_),
    .Z(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4162_ (.I(\as2650.r0[1] ),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4163_ (.I(_3698_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4164_ (.A1(_3699_),
    .A2(_3492_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4165_ (.A1(_3532_),
    .A2(_3697_),
    .B(_3700_),
    .C(_3550_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4166_ (.I(\as2650.r123_2[0][1] ),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4167_ (.I0(\as2650.r123[0][1] ),
    .I1(_3702_),
    .I2(\as2650.r123[2][1] ),
    .I3(\as2650.r123_2[2][1] ),
    .S0(_3477_),
    .S1(_3492_),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4168_ (.A1(_3520_),
    .A2(_3703_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4169_ (.A1(_3701_),
    .A2(_3704_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4170_ (.I(_3705_),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4171_ (.I(_3706_),
    .Z(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4172_ (.I(_3707_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4173_ (.A1(_3670_),
    .A2(_3696_),
    .B1(_3708_),
    .B2(_3695_),
    .C(_3642_),
    .ZN(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4174_ (.A1(_3642_),
    .A2(_3664_),
    .B(_3709_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4175_ (.I(\as2650.r0[0] ),
    .Z(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4176_ (.I(_3711_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4177_ (.I(_3712_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4178_ (.I(_3713_),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4179_ (.I(_3714_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_3631_),
    .Z(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4181_ (.A1(_3715_),
    .A2(_3716_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4182_ (.A1(_3693_),
    .A2(_3609_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4183_ (.I(_3718_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4184_ (.A1(_3637_),
    .A2(_3710_),
    .B(_3717_),
    .C(_3719_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4185_ (.I(_3592_),
    .Z(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4186_ (.A1(_3621_),
    .A2(_3721_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4187_ (.I(_3722_),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4188_ (.I(_3688_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4189_ (.I(\as2650.addr_buff[5] ),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4190_ (.A1(\as2650.addr_buff[6] ),
    .A2(_3725_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4191_ (.I(\as2650.addr_buff[6] ),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4192_ (.A1(_3727_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4193_ (.A1(_3726_),
    .A2(_3728_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4194_ (.A1(_3724_),
    .A2(_3729_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4195_ (.I(_3730_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4196_ (.A1(_3719_),
    .A2(_3731_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_3723_),
    .A2(_3732_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4198_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4199_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3734_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4200_ (.I(_3554_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4201_ (.A1(_3736_),
    .A2(_3555_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4202_ (.A1(_3735_),
    .A2(_3737_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4203_ (.A1(_3724_),
    .A2(_3738_),
    .Z(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4204_ (.I(_3739_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4205_ (.A1(_3720_),
    .A2(_3733_),
    .B1(_3740_),
    .B2(_3723_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4206_ (.I(_3715_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(\as2650.r123[0][0] ),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4208_ (.I(_3743_),
    .Z(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4209_ (.I(_3744_),
    .Z(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4210_ (.I(_3516_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4211_ (.A1(_3742_),
    .A2(_3745_),
    .A3(_3746_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4212_ (.I(_3563_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4213_ (.I(_3748_),
    .Z(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4214_ (.A1(_3517_),
    .A2(_3741_),
    .B(_3747_),
    .C(_3749_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4215_ (.A1(_3538_),
    .A2(_3562_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4216_ (.I(_3500_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_3752_),
    .Z(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4218_ (.A1(_3753_),
    .A2(_3574_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4219_ (.I(_3754_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4220_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3623_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4221_ (.I(_3683_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4222_ (.I(_3686_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4223_ (.I(\as2650.holding_reg[0] ),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4224_ (.A1(_3757_),
    .A2(_3758_),
    .B(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4225_ (.A1(_3624_),
    .A2(_3688_),
    .B(_3756_),
    .C(_3760_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4226_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3501_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4227_ (.A1(_3502_),
    .A2(_3724_),
    .B(_3760_),
    .C(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4228_ (.A1(_3761_),
    .A2(_3763_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4229_ (.I(_3764_),
    .ZN(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4230_ (.A1(_3761_),
    .A2(_3763_),
    .B(\as2650.psl[3] ),
    .C(\as2650.carry ),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4231_ (.I(\as2650.carry ),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4232_ (.A1(\as2650.psl[3] ),
    .A2(_3767_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4233_ (.A1(_3768_),
    .A2(_3764_),
    .ZN(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4234_ (.I(_3505_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4235_ (.A1(_3770_),
    .A2(_3595_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4236_ (.I(_3771_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4237_ (.A1(_3753_),
    .A2(_3772_),
    .ZN(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4238_ (.A1(_3766_),
    .A2(_3769_),
    .A3(_3773_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4239_ (.I(_3625_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4240_ (.I(_3775_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4241_ (.A1(_3776_),
    .A2(_3691_),
    .B(_3756_),
    .ZN(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4242_ (.A1(_3663_),
    .A2(_3765_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4243_ (.I(_3508_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4244_ (.A1(_3753_),
    .A2(_3779_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4245_ (.A1(_3662_),
    .A2(_3764_),
    .B(_3780_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4246_ (.I(_3752_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4247_ (.A1(_3757_),
    .A2(_3758_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4248_ (.I(_3783_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4249_ (.I(_3762_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4250_ (.A1(_3624_),
    .A2(_3784_),
    .B(_3785_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4251_ (.I(_3505_),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4252_ (.A1(_3787_),
    .A2(_3578_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4253_ (.A1(_3782_),
    .A2(_3786_),
    .B(_3788_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4254_ (.A1(_3772_),
    .A2(_3777_),
    .B1(_3778_),
    .B2(_3781_),
    .C(_3789_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4255_ (.A1(_3774_),
    .A2(_3790_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4256_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3784_),
    .ZN(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4257_ (.A1(_3782_),
    .A2(_3788_),
    .ZN(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4258_ (.A1(_3792_),
    .A2(_3793_),
    .B(_3755_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4259_ (.A1(_3755_),
    .A2(_3765_),
    .B1(_3791_),
    .B2(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4260_ (.I(_3795_),
    .Z(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4261_ (.A1(_3751_),
    .A2(_3796_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4262_ (.A1(_3750_),
    .A2(_3797_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4263_ (.I(_3798_),
    .ZN(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4264_ (.I(_3634_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4265_ (.A1(\as2650.r123[2][0] ),
    .A2(_3636_),
    .B1(_3799_),
    .B2(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4266_ (.A1(_3518_),
    .A2(_3801_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4267_ (.I(_3748_),
    .Z(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4268_ (.I(\as2650.holding_reg[1] ),
    .Z(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4269_ (.A1(_3803_),
    .A2(_3624_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4270_ (.A1(_3625_),
    .A2(_3705_),
    .B(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4271_ (.A1(_3754_),
    .A2(_3805_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4272_ (.I(_3557_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4273_ (.I(_3807_),
    .Z(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4274_ (.A1(_3770_),
    .A2(_3506_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4275_ (.A1(_3808_),
    .A2(_3809_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4276_ (.A1(_3701_),
    .A2(_3704_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4277_ (.A1(\as2650.holding_reg[1] ),
    .A2(_3811_),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4278_ (.I(_3812_),
    .Z(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4279_ (.A1(_3808_),
    .A2(_3771_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4280_ (.I(_3814_),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4281_ (.I(_3811_),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4282_ (.A1(\as2650.holding_reg[1] ),
    .A2(_3816_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4283_ (.A1(_3812_),
    .A2(_3817_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4284_ (.A1(_3760_),
    .A2(_3786_),
    .B1(_3761_),
    .B2(_3663_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4285_ (.A1(_3818_),
    .A2(_3819_),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4286_ (.A1(_3808_),
    .A2(_3779_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4287_ (.A1(_3792_),
    .A2(_3766_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4288_ (.A1(_3818_),
    .A2(_3822_),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_3752_),
    .A2(_3809_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4290_ (.A1(_3803_),
    .A2(_3549_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4291_ (.A1(_3549_),
    .A2(_3707_),
    .B(_3825_),
    .C(_3771_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4292_ (.A1(_3821_),
    .A2(_3823_),
    .B(_3824_),
    .C(_3826_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4293_ (.A1(_3815_),
    .A2(_3820_),
    .B(_3827_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4294_ (.I(_3788_),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4295_ (.A1(_3782_),
    .A2(_3817_),
    .B(_3829_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4296_ (.A1(_3810_),
    .A2(_3813_),
    .B1(_3828_),
    .B2(_3830_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4297_ (.A1(_3806_),
    .A2(_3831_),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_3832_),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4299_ (.I(_3699_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4300_ (.I(_3834_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4301_ (.I(_3835_),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4302_ (.I(\as2650.r123[0][1] ),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4303_ (.I(_3837_),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4304_ (.I(_3838_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4305_ (.A1(_3836_),
    .A2(_3714_),
    .A3(_3744_),
    .A4(_3839_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4306_ (.I(_3539_),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4307_ (.I(_3836_),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4308_ (.I(_3842_),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4309_ (.A1(_3843_),
    .A2(_3745_),
    .B1(_3839_),
    .B2(_3742_),
    .ZN(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4310_ (.A1(_3841_),
    .A2(_3844_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4311_ (.I(\as2650.addr_buff[7] ),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4312_ (.A1(_3846_),
    .A2(_3607_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4313_ (.I(_3542_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4314_ (.A1(_3848_),
    .A2(_3603_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4315_ (.A1(_3621_),
    .A2(_3847_),
    .A3(_3849_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(_3850_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4317_ (.I(_3691_),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_3620_),
    .A2(_3598_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4319_ (.I(_3853_),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4320_ (.A1(_3577_),
    .A2(_3582_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4321_ (.A1(_3619_),
    .A2(_3855_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4322_ (.I(_3856_),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4323_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123_2[1][2] ),
    .S(_3647_),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4324_ (.I(\as2650.r0[2] ),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4325_ (.I(_3859_),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4326_ (.I(_3860_),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4327_ (.A1(_3861_),
    .A2(_3614_),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4328_ (.I(_3550_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4329_ (.A1(_3532_),
    .A2(_3858_),
    .B(_3862_),
    .C(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4330_ (.I(\as2650.r123[0][2] ),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4331_ (.I(_3865_),
    .Z(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4332_ (.I(\as2650.r123_2[0][2] ),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(_3867_),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4334_ (.I0(_3866_),
    .I1(_3868_),
    .I2(\as2650.r123[2][2] ),
    .I3(\as2650.r123_2[2][2] ),
    .S0(_3478_),
    .S1(_3614_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4335_ (.A1(_3521_),
    .A2(_3869_),
    .ZN(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4336_ (.A1(_3864_),
    .A2(_3870_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4337_ (.I(_3871_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4338_ (.I(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4339_ (.I(_3873_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(_3668_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4341_ (.A1(_3557_),
    .A2(_3626_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4342_ (.A1(_3540_),
    .A2(_3876_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4343_ (.A1(_3566_),
    .A2(_3560_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(_3690_),
    .A2(_3878_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4345_ (.A1(_3877_),
    .A2(_3690_),
    .B(_3879_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4346_ (.A1(_3707_),
    .A2(_3880_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4347_ (.I(net6),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4348_ (.I(_3882_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4349_ (.I(_3668_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4350_ (.A1(_3883_),
    .A2(_3884_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4351_ (.I(_3856_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4352_ (.A1(_3875_),
    .A2(_3881_),
    .B(_3885_),
    .C(_3886_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4353_ (.I(_3853_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4354_ (.A1(_3857_),
    .A2(_3874_),
    .B(_3887_),
    .C(_3888_),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4355_ (.I(_3630_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4356_ (.A1(_3852_),
    .A2(_3854_),
    .B(_3889_),
    .C(_3890_),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4357_ (.A1(_3843_),
    .A2(_3716_),
    .B(_3851_),
    .C(_3891_),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4358_ (.A1(_3687_),
    .A2(_3705_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4359_ (.I(_3893_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4360_ (.I(_3726_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4361_ (.A1(\as2650.addr_buff[6] ),
    .A2(_3725_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4362_ (.A1(_3724_),
    .A2(_3895_),
    .B(_3896_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4363_ (.A1(_3894_),
    .A2(_3897_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4364_ (.A1(_3894_),
    .A2(_3897_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_3898_),
    .A2(_3899_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4366_ (.A1(_3621_),
    .A2(_3721_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4367_ (.A1(_3719_),
    .A2(_3900_),
    .B(_3901_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4368_ (.I(_3735_),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4369_ (.A1(_3554_),
    .A2(_3734_),
    .ZN(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4370_ (.A1(_3688_),
    .A2(_3903_),
    .B(_3904_),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4371_ (.A1(_3894_),
    .A2(_3905_),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4372_ (.A1(_3894_),
    .A2(_3905_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4373_ (.A1(_3906_),
    .A2(_3907_),
    .Z(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4374_ (.I(_3901_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4375_ (.A1(_3892_),
    .A2(_3902_),
    .B1(_3908_),
    .B2(_3909_),
    .C(_3516_),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4376_ (.A1(_3840_),
    .A2(_3845_),
    .B(_3910_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4377_ (.A1(_3749_),
    .A2(_3911_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4378_ (.A1(_3802_),
    .A2(_3833_),
    .B(_3912_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4379_ (.I(_3913_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4380_ (.A1(\as2650.r123[2][1] ),
    .A2(_3636_),
    .B1(_3914_),
    .B2(_3800_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4381_ (.A1(_3518_),
    .A2(_3915_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(_3809_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4383_ (.I(\as2650.holding_reg[2] ),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4384_ (.A1(_3917_),
    .A2(_3874_),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4385_ (.I(_3773_),
    .Z(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4386_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3872_),
    .Z(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4387_ (.I(_3920_),
    .Z(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4388_ (.A1(_3812_),
    .A2(_3817_),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4389_ (.A1(_3792_),
    .A2(_3766_),
    .B(_3922_),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4390_ (.A1(_3813_),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4391_ (.A1(_3921_),
    .A2(_3924_),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4392_ (.A1(_3803_),
    .A2(_3816_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4393_ (.A1(_3805_),
    .A2(_3926_),
    .B1(_3922_),
    .B2(_3819_),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4394_ (.A1(_3921_),
    .A2(_3927_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4395_ (.A1(_3864_),
    .A2(_3870_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4396_ (.I(_3929_),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4397_ (.A1(_3917_),
    .A2(_3775_),
    .ZN(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4398_ (.A1(_3776_),
    .A2(_3930_),
    .B(_3931_),
    .C(_3814_),
    .ZN(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4399_ (.A1(_3815_),
    .A2(_3928_),
    .B(_3932_),
    .C(_3773_),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4400_ (.I(_3808_),
    .Z(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4401_ (.A1(_3934_),
    .A2(_3788_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4402_ (.A1(_3919_),
    .A2(_3925_),
    .B(_3933_),
    .C(_3935_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4403_ (.I(_3793_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4404_ (.A1(_3916_),
    .A2(_3918_),
    .B(_3936_),
    .C(_3937_),
    .ZN(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4405_ (.I(_3810_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4406_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3872_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4407_ (.A1(_3782_),
    .A2(_3574_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4408_ (.A1(_3939_),
    .A2(_0261_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_3755_),
    .A2(_3921_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4410_ (.A1(_3938_),
    .A2(_0263_),
    .B(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4411_ (.I(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4412_ (.I(_3516_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4413_ (.A1(_3689_),
    .A2(_3705_),
    .B(_3929_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4414_ (.A1(_3784_),
    .A2(_3811_),
    .A3(_3871_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4415_ (.A1(_3904_),
    .A2(_0268_),
    .A3(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4416_ (.A1(_3736_),
    .A2(_3555_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4417_ (.A1(_0271_),
    .A2(_3904_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4418_ (.A1(_3757_),
    .A2(_3758_),
    .B1(_3701_),
    .B2(_3704_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4419_ (.A1(_3872_),
    .A2(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4420_ (.I(_0271_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4421_ (.A1(_0272_),
    .A2(_3873_),
    .B1(_0274_),
    .B2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4422_ (.A1(_0270_),
    .A2(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4423_ (.I(_3861_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4424_ (.I(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4425_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4426_ (.I(_3718_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4427_ (.A1(_3689_),
    .A2(_3706_),
    .A3(_3878_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4428_ (.A1(_3877_),
    .A2(_3690_),
    .A3(_3706_),
    .B(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4429_ (.A1(_3873_),
    .A2(_0283_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4430_ (.I(net7),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_0285_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4432_ (.I(_0286_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4433_ (.I(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4434_ (.I(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4435_ (.A1(_0289_),
    .A2(_3678_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4436_ (.A1(_3678_),
    .A2(_0284_),
    .B(_0290_),
    .C(_3694_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4437_ (.A1(_3479_),
    .A2(\as2650.r123[1][3] ),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4438_ (.A1(_3648_),
    .A2(\as2650.r123_2[1][3] ),
    .B(_3493_),
    .C(_3863_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4439_ (.I(\as2650.r0[3] ),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4440_ (.I(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4442_ (.A1(_0296_),
    .A2(_3615_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(\as2650.r123[0][3] ),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4444_ (.I(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4445_ (.I0(_0299_),
    .I1(\as2650.r123_2[0][3] ),
    .I2(\as2650.r123[2][3] ),
    .I3(\as2650.r123_2[2][3] ),
    .S0(_3478_),
    .S1(_3492_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_3520_),
    .A2(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4447_ (.A1(_0292_),
    .A2(_0293_),
    .B(_0297_),
    .C(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4448_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4449_ (.I(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4450_ (.I(_0304_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4451_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4452_ (.I(_0306_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4453_ (.A1(_3857_),
    .A2(_0307_),
    .B(_3888_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4454_ (.A1(_3854_),
    .A2(_3708_),
    .B1(_0291_),
    .B2(_0308_),
    .C(_3631_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4455_ (.A1(_0280_),
    .A2(_3716_),
    .B(_0281_),
    .C(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4456_ (.I(_3585_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4457_ (.I(_0311_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4458_ (.A1(_3600_),
    .A2(_3607_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4459_ (.I(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4460_ (.I(_3603_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4461_ (.A1(_0312_),
    .A2(_3693_),
    .A3(_0314_),
    .A4(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4462_ (.A1(_3896_),
    .A2(_0268_),
    .A3(_0269_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4463_ (.I(_3729_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4464_ (.A1(_3727_),
    .A2(_3606_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4465_ (.A1(_0318_),
    .A2(_3873_),
    .B1(_0274_),
    .B2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4466_ (.A1(_0317_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4467_ (.A1(_0316_),
    .A2(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4468_ (.A1(_3722_),
    .A2(_0310_),
    .A3(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4469_ (.A1(_3723_),
    .A2(_0277_),
    .B(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4470_ (.A1(_3681_),
    .A2(\as2650.r123[0][2] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4471_ (.A1(_3836_),
    .A2(_3838_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(_3861_),
    .A2(_3743_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4473_ (.A1(_0278_),
    .A2(_3835_),
    .A3(_3744_),
    .A4(_3838_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4474_ (.A1(_0326_),
    .A2(_0327_),
    .B(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4475_ (.A1(_0325_),
    .A2(_0329_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4476_ (.A1(_3840_),
    .A2(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4477_ (.A1(_3746_),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4478_ (.I(_3748_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4479_ (.A1(_0267_),
    .A2(_0324_),
    .B(_0332_),
    .C(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4480_ (.A1(_3802_),
    .A2(_0266_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4481_ (.I(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4482_ (.A1(\as2650.r123[2][2] ),
    .A2(_3636_),
    .B1(_0336_),
    .B2(_3800_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4483_ (.A1(_3518_),
    .A2(_0337_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4484_ (.I(_0262_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4485_ (.I(\as2650.holding_reg[3] ),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4486_ (.I(_0303_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4487_ (.A1(_0339_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4488_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0304_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4489_ (.I(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4490_ (.A1(_0341_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4491_ (.I(_0341_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4492_ (.A1(_0345_),
    .A2(_0343_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4493_ (.I(_3864_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4494_ (.I(_3870_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _4495_ (.A1(_3917_),
    .A2(_0347_),
    .A3(_0348_),
    .B1(_3813_),
    .B2(_3923_),
    .B3(_0261_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4496_ (.A1(_0346_),
    .A2(_0349_),
    .B(_3919_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4497_ (.A1(_0346_),
    .A2(_0349_),
    .B(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4498_ (.A1(_3502_),
    .A2(_3930_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4499_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3503_),
    .B(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4500_ (.A1(_3920_),
    .A2(_3927_),
    .B1(_0353_),
    .B2(_0261_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4501_ (.A1(_0344_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(_3776_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(_0356_),
    .A2(_0305_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4504_ (.I(_3503_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4505_ (.I(_0358_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4506_ (.A1(_0339_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4507_ (.A1(_3772_),
    .A2(_0357_),
    .A3(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4508_ (.A1(_3780_),
    .A2(_0355_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4509_ (.I0(_0339_),
    .I1(_0340_),
    .S(_3502_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4510_ (.A1(_3934_),
    .A2(_0363_),
    .B(_3916_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4511_ (.A1(_0351_),
    .A2(_0362_),
    .B(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4512_ (.A1(_3937_),
    .A2(_0345_),
    .B(_3755_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4513_ (.A1(_0365_),
    .A2(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4514_ (.A1(_0338_),
    .A2(_0344_),
    .B(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4515_ (.I(_3901_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _4516_ (.A1(_3757_),
    .A2(_3758_),
    .B1(_3701_),
    .B2(_3704_),
    .C1(_3864_),
    .C2(_3870_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4517_ (.A1(_0370_),
    .A2(_0303_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4518_ (.I(_3737_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _4519_ (.A1(_0269_),
    .A2(_0304_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4520_ (.A1(_0272_),
    .A2(_0340_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4521_ (.A1(_0372_),
    .A2(_0373_),
    .B(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4522_ (.A1(_0275_),
    .A2(_0371_),
    .B(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4523_ (.I(_3728_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4524_ (.A1(_0318_),
    .A2(_0305_),
    .B1(_0371_),
    .B2(_0319_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4525_ (.A1(_0377_),
    .A2(_0373_),
    .B(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4526_ (.I(_0379_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4527_ (.A1(_3498_),
    .A2(_3876_),
    .A3(_0370_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4528_ (.A1(_3689_),
    .A2(_3706_),
    .A3(_3878_),
    .A4(_3930_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_0381_),
    .A2(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4530_ (.A1(_0305_),
    .A2(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4531_ (.A1(_3678_),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4532_ (.I(net8),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4533_ (.I(_0386_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4535_ (.A1(_0388_),
    .A2(_3669_),
    .B(_3694_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(\as2650.r0[4] ),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4538_ (.I(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4539_ (.I(\as2650.r123[0][4] ),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4540_ (.I(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4541_ (.I0(_0394_),
    .I1(\as2650.r123_2[0][4] ),
    .I2(\as2650.r123[2][4] ),
    .I3(\as2650.r123_2[2][4] ),
    .S0(_3647_),
    .S1(_3493_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4542_ (.I(_3478_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4543_ (.A1(_0396_),
    .A2(\as2650.r123[1][4] ),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4544_ (.A1(_3649_),
    .A2(\as2650.r123_2[1][4] ),
    .B(_3494_),
    .C(_3863_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4545_ (.A1(_0397_),
    .A2(_0398_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4546_ (.A1(_0392_),
    .A2(_3617_),
    .B1(_0395_),
    .B2(_3522_),
    .C(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4547_ (.I(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_0401_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(_3641_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4550_ (.A1(_0385_),
    .A2(_0389_),
    .B1(_0402_),
    .B2(_3695_),
    .C(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4551_ (.A1(_3642_),
    .A2(_3874_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4552_ (.I(_0296_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4553_ (.I(_0406_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4554_ (.A1(_0407_),
    .A2(_3632_),
    .B(_3850_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4555_ (.A1(_3637_),
    .A2(_0405_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4556_ (.A1(_0316_),
    .A2(_0380_),
    .B(_0409_),
    .C(_3909_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4557_ (.A1(_0369_),
    .A2(_0376_),
    .B(_0410_),
    .C(_0267_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4558_ (.I(_3539_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4559_ (.A1(_3840_),
    .A2(_0330_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4560_ (.A1(_0326_),
    .A2(_0327_),
    .B(_0328_),
    .C(_0325_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(\as2650.r0[1] ),
    .A2(_0298_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4562_ (.A1(_0325_),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4563_ (.A1(_3834_),
    .A2(_3866_),
    .B1(_0299_),
    .B2(_3712_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4564_ (.A1(_0416_),
    .A2(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4565_ (.A1(_0296_),
    .A2(_3743_),
    .B1(_3837_),
    .B2(_3861_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4566_ (.A1(_0295_),
    .A2(\as2650.r123[0][1] ),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4567_ (.A1(_0327_),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4568_ (.A1(_0419_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4569_ (.A1(_0418_),
    .A2(_0422_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4570_ (.A1(_0328_),
    .A2(_0414_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4571_ (.A1(_0328_),
    .A2(_0414_),
    .A3(_0423_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4572_ (.A1(_0424_),
    .A2(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4573_ (.A1(_0413_),
    .A2(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4574_ (.A1(_0413_),
    .A2(_0426_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4575_ (.A1(_0412_),
    .A2(_0427_),
    .A3(_0428_),
    .B(_0333_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4576_ (.A1(_3749_),
    .A2(_0368_),
    .B1(_0411_),
    .B2(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4577_ (.I(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4578_ (.A1(\as2650.r123[2][3] ),
    .A2(_3636_),
    .B1(_0431_),
    .B2(_3800_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4579_ (.A1(_3518_),
    .A2(_0432_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_3635_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4581_ (.I(_3754_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4582_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4583_ (.I(_3815_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_0391_),
    .A2(_3616_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4585_ (.A1(_3521_),
    .A2(_0395_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4586_ (.A1(_0397_),
    .A2(_0398_),
    .B(_0437_),
    .C(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4587_ (.I(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4589_ (.I(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4590_ (.I(\as2650.holding_reg[4] ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4591_ (.A1(_0443_),
    .A2(_0401_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4592_ (.A1(_0442_),
    .A2(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4593_ (.A1(_0341_),
    .A2(_0363_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4594_ (.A1(_0344_),
    .A2(_0354_),
    .B(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4595_ (.A1(_0445_),
    .A2(_0447_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4596_ (.I(_0440_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4597_ (.A1(_0443_),
    .A2(_0356_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4598_ (.A1(_0356_),
    .A2(_0449_),
    .B(_0450_),
    .C(_0436_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4599_ (.A1(_0436_),
    .A2(_0448_),
    .B(_0451_),
    .C(_3919_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4600_ (.I(_3821_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4601_ (.A1(_0342_),
    .A2(_0349_),
    .B(_0345_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4602_ (.A1(_0445_),
    .A2(_0454_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4603_ (.A1(\as2650.holding_reg[4] ),
    .A2(_3625_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4604_ (.A1(_0358_),
    .A2(_0440_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4605_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_3916_),
    .A2(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4607_ (.A1(_0453_),
    .A2(_0455_),
    .B(_0459_),
    .C(_3939_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4608_ (.A1(_3937_),
    .A2(_0442_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4609_ (.A1(_0452_),
    .A2(_0460_),
    .B(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4610_ (.A1(_0441_),
    .A2(_0444_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_0434_),
    .A2(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4612_ (.A1(_0435_),
    .A2(_0462_),
    .B(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4613_ (.A1(_0416_),
    .A2(_0420_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_0391_),
    .A2(\as2650.r123[0][0] ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4615_ (.A1(_0466_),
    .A2(_0467_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4616_ (.A1(_3681_),
    .A2(_0393_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4617_ (.A1(_0415_),
    .A2(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(_0415_),
    .A2(_0469_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_0470_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4620_ (.A1(_3860_),
    .A2(_3865_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4621_ (.A1(_0472_),
    .A2(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4622_ (.A1(_0468_),
    .A2(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4623_ (.A1(_0418_),
    .A2(_0422_),
    .B(_0421_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4624_ (.A1(_0475_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4625_ (.A1(_0424_),
    .A2(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4626_ (.A1(_0428_),
    .A2(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(_0428_),
    .A2(_0478_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4628_ (.A1(_3746_),
    .A2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4629_ (.A1(_3783_),
    .A2(_3811_),
    .A3(_3871_),
    .A4(_0302_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4630_ (.A1(_0439_),
    .A2(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4631_ (.A1(_0370_),
    .A2(_0303_),
    .A3(_0439_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4632_ (.I(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4633_ (.A1(_0370_),
    .A2(_0304_),
    .B(_0439_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4634_ (.A1(_0485_),
    .A2(_0486_),
    .B(_3895_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4635_ (.I(_3729_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(_0488_),
    .A2(_0401_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4637_ (.A1(_3896_),
    .A2(_0483_),
    .B(_0487_),
    .C(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4638_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4639_ (.I(_0392_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4640_ (.I0(_0382_),
    .I1(_0381_),
    .S(_0340_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4641_ (.A1(_0440_),
    .A2(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4642_ (.I(net9),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(_0495_),
    .A2(_3884_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4644_ (.A1(_3875_),
    .A2(_0494_),
    .B(_0496_),
    .C(_3886_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4645_ (.I(\as2650.r0[5] ),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4646_ (.I(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(\as2650.r123[0][5] ),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(\as2650.r123_2[0][5] ),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4649_ (.I0(_0500_),
    .I1(_0501_),
    .I2(\as2650.r123[2][5] ),
    .I3(\as2650.r123_2[2][5] ),
    .S0(_3479_),
    .S1(_3494_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4650_ (.A1(_0396_),
    .A2(\as2650.r123[1][5] ),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4651_ (.A1(_3649_),
    .A2(\as2650.r123_2[1][5] ),
    .B(_3494_),
    .C(_3551_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4652_ (.A1(_0503_),
    .A2(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4653_ (.A1(_0499_),
    .A2(_3617_),
    .B1(_0502_),
    .B2(_3522_),
    .C(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4654_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4655_ (.A1(_3694_),
    .A2(_0507_),
    .B(_0403_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4656_ (.A1(_0403_),
    .A2(_0306_),
    .B1(_0497_),
    .B2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4657_ (.A1(_3890_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4658_ (.A1(_0492_),
    .A2(_3632_),
    .B(_3850_),
    .C(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4659_ (.A1(_0281_),
    .A2(_0491_),
    .B(_0511_),
    .C(_3722_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4660_ (.A1(_0485_),
    .A2(_0486_),
    .B(_3903_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4661_ (.I(_3738_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_0514_),
    .A2(_0401_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4663_ (.A1(_3904_),
    .A2(_0483_),
    .B(_0513_),
    .C(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4664_ (.I(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4665_ (.A1(_3909_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4666_ (.A1(_0412_),
    .A2(_0512_),
    .A3(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4667_ (.A1(_0479_),
    .A2(_0481_),
    .B(_0519_),
    .C(_0333_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4668_ (.A1(_3802_),
    .A2(_0465_),
    .B(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4669_ (.I(_0521_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4670_ (.A1(\as2650.r123[2][4] ),
    .A2(_0433_),
    .B1(_0522_),
    .B2(_3634_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4671_ (.A1(_3517_),
    .A2(_0523_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4672_ (.I(_3841_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4673_ (.I(_3634_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_0499_),
    .A2(_3616_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4675_ (.A1(_3522_),
    .A2(_0502_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4676_ (.A1(_0503_),
    .A2(_0504_),
    .B(_0526_),
    .C(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4677_ (.I(_0528_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4678_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(\as2650.holding_reg[5] ),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4680_ (.I(_0529_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4681_ (.A1(_0531_),
    .A2(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(_0530_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4683_ (.A1(_0530_),
    .A2(_0533_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(_0442_),
    .A2(_0458_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4685_ (.A1(_0463_),
    .A2(_0447_),
    .B(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4686_ (.A1(_0535_),
    .A2(_0537_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4687_ (.I(_0359_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4688_ (.A1(_0539_),
    .A2(_0507_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4689_ (.A1(_0531_),
    .A2(_0539_),
    .B(_0436_),
    .C(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4690_ (.A1(_0436_),
    .A2(_0538_),
    .B(_0541_),
    .C(_3919_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4691_ (.A1(_0342_),
    .A2(_0349_),
    .B(_0442_),
    .C(_0345_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4692_ (.A1(_0444_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4693_ (.A1(_0535_),
    .A2(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_0453_),
    .A2(_0545_),
    .B(_3824_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4695_ (.I(_3753_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4696_ (.A1(_0547_),
    .A2(_0530_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4697_ (.A1(_0542_),
    .A2(_0546_),
    .B1(_0548_),
    .B2(_3829_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4698_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0532_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4699_ (.A1(_3937_),
    .A2(_0550_),
    .B(_0434_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4700_ (.A1(_0435_),
    .A2(_0534_),
    .B1(_0549_),
    .B2(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4701_ (.I(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4702_ (.A1(_0400_),
    .A2(_0482_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4703_ (.A1(_0529_),
    .A2(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4704_ (.A1(_0528_),
    .A2(_0485_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4705_ (.A1(_0275_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4706_ (.A1(_0514_),
    .A2(_0506_),
    .B1(_0555_),
    .B2(_0372_),
    .C(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4707_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4708_ (.I(_0499_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4709_ (.I(_0402_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4710_ (.A1(_0396_),
    .A2(\as2650.r123[1][6] ),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4711_ (.A1(_3649_),
    .A2(\as2650.r123_2[1][6] ),
    .B(_3493_),
    .C(_3863_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4712_ (.I(\as2650.r0[6] ),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4713_ (.A1(_0564_),
    .A2(_3616_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _4714_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .I2(\as2650.r123[2][6] ),
    .I3(\as2650.r123_2[2][6] ),
    .S0(_3647_),
    .S1(_3614_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4715_ (.A1(_3521_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4716_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0565_),
    .C(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4717_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4718_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4719_ (.A1(_3541_),
    .A2(_3876_),
    .A3(_0485_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4720_ (.A1(_3807_),
    .A2(_3626_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4721_ (.A1(_3498_),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4722_ (.A1(_0573_),
    .A2(_0554_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4723_ (.A1(_0571_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4724_ (.A1(_0532_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4725_ (.I(net1),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4726_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4727_ (.I(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4728_ (.I(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4729_ (.A1(_0580_),
    .A2(_3884_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4730_ (.A1(_3669_),
    .A2(_0576_),
    .B(_0581_),
    .C(_3886_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4731_ (.A1(_3857_),
    .A2(_0570_),
    .B(_0582_),
    .C(_3888_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4732_ (.A1(_3854_),
    .A2(_0561_),
    .B(_0583_),
    .C(_3890_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4733_ (.A1(_0560_),
    .A2(_3637_),
    .B(_3851_),
    .C(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4734_ (.A1(_0319_),
    .A2(_0556_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4735_ (.A1(_0488_),
    .A2(_0507_),
    .B1(_0555_),
    .B2(_0377_),
    .C(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4736_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4737_ (.A1(_0316_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4738_ (.A1(_0585_),
    .A2(_0589_),
    .B(_0369_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4739_ (.A1(_0369_),
    .A2(_0559_),
    .B(_0590_),
    .C(_0267_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4740_ (.A1(_0424_),
    .A2(_0477_),
    .B(_0480_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4741_ (.A1(_0475_),
    .A2(_0476_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4742_ (.I(_0474_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(_0468_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4744_ (.A1(_0406_),
    .A2(_3838_),
    .A3(_0416_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4745_ (.A1(_0466_),
    .A2(_0467_),
    .B(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4746_ (.A1(_3711_),
    .A2(_0500_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4747_ (.A1(_3860_),
    .A2(_3698_),
    .A3(_0298_),
    .A4(_0393_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4748_ (.A1(_3860_),
    .A2(_0298_),
    .B1(_0394_),
    .B2(_3698_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4749_ (.A1(_0599_),
    .A2(_0600_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_0295_),
    .A2(_3865_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4751_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4752_ (.A1(_0598_),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4753_ (.A1(_0472_),
    .A2(_0473_),
    .B(_0470_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4754_ (.A1(_0391_),
    .A2(_3837_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4755_ (.A1(_0605_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4756_ (.A1(_0498_),
    .A2(_3743_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4757_ (.A1(_0607_),
    .A2(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4758_ (.A1(_0604_),
    .A2(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4759_ (.A1(_0595_),
    .A2(_0597_),
    .A3(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4760_ (.A1(_0593_),
    .A2(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4761_ (.A1(_0592_),
    .A2(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4762_ (.A1(_0524_),
    .A2(_0613_),
    .B(_0333_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4763_ (.A1(_0591_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4764_ (.A1(_3751_),
    .A2(_0553_),
    .B(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4765_ (.A1(\as2650.r123[2][5] ),
    .A2(_0433_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4766_ (.A1(_0525_),
    .A2(_0616_),
    .B(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4767_ (.A1(_0524_),
    .A2(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4768_ (.I(_0619_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4769_ (.A1(_0593_),
    .A2(_0611_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4770_ (.A1(_0592_),
    .A2(_0612_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4771_ (.A1(_0604_),
    .A2(_0609_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4772_ (.I(_0606_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4773_ (.A1(_0607_),
    .A2(_0608_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4774_ (.A1(_0605_),
    .A2(_0623_),
    .B(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_0598_),
    .A2(_0603_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4776_ (.A1(_0294_),
    .A2(\as2650.r123[0][3] ),
    .B1(_0393_),
    .B2(_3859_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4777_ (.A1(_0294_),
    .A2(_3859_),
    .A3(\as2650.r123[0][3] ),
    .A4(\as2650.r123[0][4] ),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4778_ (.A1(_0627_),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(_0390_),
    .A2(_3865_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4780_ (.A1(_0629_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4781_ (.A1(_3711_),
    .A2(\as2650.r123[0][6] ),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4782_ (.A1(_3698_),
    .A2(\as2650.r123[0][5] ),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4783_ (.A1(_0632_),
    .A2(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4784_ (.A1(_0631_),
    .A2(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4785_ (.A1(_0626_),
    .A2(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4786_ (.I(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4787_ (.A1(_0601_),
    .A2(_0602_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4788_ (.A1(_0599_),
    .A2(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4789_ (.A1(_0499_),
    .A2(_3837_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_0564_),
    .A2(_3744_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4791_ (.A1(_0639_),
    .A2(_0640_),
    .A3(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4792_ (.A1(_0637_),
    .A2(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4793_ (.A1(_0622_),
    .A2(_0625_),
    .A3(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4794_ (.A1(_0595_),
    .A2(_0610_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4795_ (.A1(_0595_),
    .A2(_0610_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4796_ (.A1(_0597_),
    .A2(_0645_),
    .B(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4797_ (.A1(_0644_),
    .A2(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4798_ (.A1(_0620_),
    .A2(_0621_),
    .A3(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4799_ (.A1(_0620_),
    .A2(_0621_),
    .B(_0648_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_0267_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4801_ (.A1(_0562_),
    .A2(_0563_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4802_ (.A1(_0564_),
    .A2(_3618_),
    .B1(_0566_),
    .B2(_3523_),
    .C(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4803_ (.A1(_0528_),
    .A2(_0484_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4804_ (.A1(_0569_),
    .A2(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4805_ (.A1(_0400_),
    .A2(_0482_),
    .A3(_0506_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4806_ (.A1(_0569_),
    .A2(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4807_ (.A1(_3737_),
    .A2(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4808_ (.A1(_0514_),
    .A2(_0653_),
    .B1(_0655_),
    .B2(_3903_),
    .C(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4809_ (.I(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4810_ (.I(_0564_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4811_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4812_ (.I(_0532_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4813_ (.I(_0653_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4814_ (.A1(_0529_),
    .A2(_0571_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4815_ (.A1(_0573_),
    .A2(_0656_),
    .B(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4816_ (.A1(_0664_),
    .A2(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4817_ (.I(net2),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4819_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4820_ (.A1(_0670_),
    .A2(_3875_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4821_ (.A1(_3669_),
    .A2(_0667_),
    .B(_0671_),
    .C(_3886_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4822_ (.A1(_3695_),
    .A2(_3660_),
    .B(_0403_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4823_ (.A1(_3642_),
    .A2(_0663_),
    .B1(_0672_),
    .B2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4824_ (.A1(_3632_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4825_ (.A1(_0662_),
    .A2(_3637_),
    .B(_3851_),
    .C(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4826_ (.A1(_3895_),
    .A2(_0655_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4827_ (.A1(_0488_),
    .A2(_0664_),
    .B1(_0657_),
    .B2(_0377_),
    .C(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4828_ (.I(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4829_ (.A1(_0316_),
    .A2(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4830_ (.A1(_3722_),
    .A2(_0676_),
    .A3(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4831_ (.A1(_3723_),
    .A2(_0660_),
    .B(_0681_),
    .C(_0412_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4832_ (.A1(_0649_),
    .A2(_0651_),
    .B(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4833_ (.I(\as2650.holding_reg[6] ),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4834_ (.A1(_0684_),
    .A2(_0664_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4835_ (.A1(_0444_),
    .A2(_0530_),
    .A3(_0543_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4836_ (.A1(_0533_),
    .A2(_0685_),
    .A3(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4837_ (.A1(_0533_),
    .A2(_0686_),
    .B(_0685_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4838_ (.A1(_3821_),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4839_ (.A1(_0687_),
    .A2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(_3780_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4841_ (.A1(_0684_),
    .A2(_0569_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4842_ (.A1(_0358_),
    .A2(_0506_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4843_ (.A1(_0531_),
    .A2(_3549_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4844_ (.A1(_0550_),
    .A2(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4845_ (.A1(_0534_),
    .A2(_0537_),
    .B(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4846_ (.A1(_0692_),
    .A2(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4847_ (.I(_0539_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4848_ (.I(_0653_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(_0684_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4850_ (.A1(_0700_),
    .A2(_0539_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4851_ (.A1(_0698_),
    .A2(_0699_),
    .B(_0701_),
    .C(_0691_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4852_ (.A1(_0691_),
    .A2(_0697_),
    .B(_0702_),
    .C(_0453_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4853_ (.A1(_0690_),
    .A2(_0703_),
    .B(_3916_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4854_ (.A1(_0684_),
    .A2(_0570_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4855_ (.I(_0570_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4856_ (.I(_3578_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4857_ (.A1(_0700_),
    .A2(_0706_),
    .B(_0547_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4858_ (.A1(_3939_),
    .A2(_0705_),
    .B(_0708_),
    .C(_0338_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4859_ (.A1(_0435_),
    .A2(_0685_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4860_ (.A1(_0704_),
    .A2(_0709_),
    .B(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4861_ (.A1(_3749_),
    .A2(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4862_ (.A1(_3802_),
    .A2(_0683_),
    .B(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4863_ (.A1(\as2650.r123[2][6] ),
    .A2(_0433_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4864_ (.A1(_0525_),
    .A2(_0713_),
    .B(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4865_ (.A1(_0524_),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(_0716_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(\as2650.holding_reg[7] ),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4868_ (.A1(_0717_),
    .A2(_3660_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4869_ (.I(_3658_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4870_ (.I(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4871_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4872_ (.A1(\as2650.holding_reg[6] ),
    .A2(_3775_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4873_ (.A1(_3775_),
    .A2(_0699_),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(_0705_),
    .A2(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4875_ (.A1(_0692_),
    .A2(_0696_),
    .B(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4876_ (.A1(_0721_),
    .A2(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4877_ (.I(_3776_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4878_ (.A1(_0356_),
    .A2(_3660_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4879_ (.A1(_0717_),
    .A2(_0727_),
    .B(_0691_),
    .C(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4880_ (.A1(_0691_),
    .A2(_0726_),
    .B(_0729_),
    .C(_0453_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4881_ (.I(_0721_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4882_ (.A1(_0700_),
    .A2(_0570_),
    .B(_0688_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4883_ (.A1(_0721_),
    .A2(_0732_),
    .B(_3821_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4884_ (.A1(_0731_),
    .A2(_0732_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4885_ (.A1(_3829_),
    .A2(_0730_),
    .A3(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_0717_),
    .A2(_0720_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4887_ (.I(_0717_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4888_ (.A1(_0737_),
    .A2(_0720_),
    .B(_3935_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4889_ (.A1(_3939_),
    .A2(_0736_),
    .B(_0738_),
    .C(_0262_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4890_ (.I(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4891_ (.A1(_0435_),
    .A2(_0718_),
    .B1(_0735_),
    .B2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4892_ (.A1(_0639_),
    .A2(_0640_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4893_ (.A1(_0639_),
    .A2(_0640_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4894_ (.A1(_0742_),
    .A2(_0641_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4895_ (.A1(_0560_),
    .A2(_3866_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4896_ (.A1(_3842_),
    .A2(\as2650.r123[0][6] ),
    .A3(_0598_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4897_ (.A1(_0279_),
    .A2(_0500_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4898_ (.A1(_0392_),
    .A2(_0299_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4899_ (.A1(_3714_),
    .A2(\as2650.r123[0][7] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4900_ (.A1(_0747_),
    .A2(_0748_),
    .A3(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4901_ (.A1(_0746_),
    .A2(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4902_ (.A1(_0744_),
    .A2(_0745_),
    .A3(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4903_ (.A1(_0644_),
    .A2(_0647_),
    .B(_0650_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_0631_),
    .A2(_0634_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4905_ (.A1(_0406_),
    .A2(_0394_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4906_ (.A1(_0627_),
    .A2(_0628_),
    .A3(_0630_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4907_ (.A1(_0628_),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4908_ (.A1(_0661_),
    .A2(_3839_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4909_ (.A1(_0755_),
    .A2(_0757_),
    .A3(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4910_ (.A1(_0622_),
    .A2(_0643_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4911_ (.A1(_0622_),
    .A2(_0643_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4912_ (.A1(_0625_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4913_ (.A1(_0598_),
    .A2(_0603_),
    .A3(_0635_),
    .B1(_0637_),
    .B2(_0642_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_3645_),
    .A2(_3745_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4915_ (.A1(_0762_),
    .A2(_0763_),
    .A3(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4916_ (.A1(_0754_),
    .A2(_0759_),
    .A3(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4917_ (.A1(_0752_),
    .A2(_0753_),
    .A3(_0766_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4918_ (.A1(_0528_),
    .A2(_0568_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4919_ (.A1(_0400_),
    .A2(_0482_),
    .A3(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4920_ (.A1(_0719_),
    .A2(_0769_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4921_ (.A1(_0653_),
    .A2(_0654_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4922_ (.A1(_3659_),
    .A2(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4923_ (.A1(_3659_),
    .A2(_0514_),
    .B1(_0770_),
    .B2(_0372_),
    .C1(_0772_),
    .C2(_3903_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4924_ (.I(_0773_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_0699_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4926_ (.A1(_3643_),
    .A2(_3691_),
    .B(_3663_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4927_ (.A1(_3877_),
    .A2(_0664_),
    .A3(_0654_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4928_ (.A1(_0719_),
    .A2(_0573_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4929_ (.A1(_0573_),
    .A2(_0770_),
    .B(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4930_ (.A1(_0777_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(net3),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4932_ (.I(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4933_ (.A1(_0782_),
    .A2(_3884_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4934_ (.A1(_3875_),
    .A2(_0780_),
    .B(_0783_),
    .C(_3856_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4935_ (.A1(_3857_),
    .A2(_0776_),
    .B(_0784_),
    .C(_3888_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4936_ (.A1(_3854_),
    .A2(_0775_),
    .B(_0785_),
    .C(_3890_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4937_ (.A1(_3645_),
    .A2(_3716_),
    .B(_3851_),
    .C(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4938_ (.A1(_0377_),
    .A2(_0770_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4939_ (.A1(_3659_),
    .A2(_0488_),
    .B1(_0772_),
    .B2(_3895_),
    .C(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4940_ (.I(_0789_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4941_ (.A1(_3719_),
    .A2(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4942_ (.A1(_0787_),
    .A2(_0791_),
    .B(_3909_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4943_ (.A1(_0369_),
    .A2(_0774_),
    .B(_0792_),
    .C(_3746_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4944_ (.A1(_3517_),
    .A2(_0767_),
    .B(_0793_),
    .C(_3751_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4945_ (.A1(_3751_),
    .A2(_0741_),
    .B(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4946_ (.A1(\as2650.r123[2][7] ),
    .A2(_0433_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4947_ (.A1(_0525_),
    .A2(_0795_),
    .B(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4948_ (.A1(_0524_),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4949_ (.I(_0798_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4950_ (.I(_3629_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4951_ (.A1(_3584_),
    .A2(_3610_),
    .A3(_0799_),
    .A4(_3613_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4952_ (.A1(_3693_),
    .A2(_0800_),
    .B(_3748_),
    .C(_3841_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4953_ (.I(_3523_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4954_ (.I(_0802_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4955_ (.A1(_0803_),
    .A2(_3534_),
    .B(_3841_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4956_ (.A1(_0801_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4957_ (.I(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_3513_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4959_ (.A1(_0807_),
    .A2(_0805_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4960_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4961_ (.A1(\as2650.r123[1][0] ),
    .A2(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4962_ (.A1(_3798_),
    .A2(_0806_),
    .B(_0810_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4963_ (.A1(\as2650.r123[1][1] ),
    .A2(_0809_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4964_ (.A1(_3913_),
    .A2(_0806_),
    .B(_0811_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4965_ (.A1(\as2650.r123[1][2] ),
    .A2(_0809_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4966_ (.A1(_0335_),
    .A2(_0806_),
    .B(_0812_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4967_ (.A1(\as2650.r123[1][3] ),
    .A2(_0809_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4968_ (.A1(_0430_),
    .A2(_0806_),
    .B(_0813_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4969_ (.I(_0805_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4970_ (.I(_0808_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4971_ (.A1(\as2650.r123[1][4] ),
    .A2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4972_ (.A1(_0521_),
    .A2(_0814_),
    .B(_0816_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(\as2650.r123[1][5] ),
    .A2(_0815_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4974_ (.A1(_0616_),
    .A2(_0814_),
    .B(_0817_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4975_ (.A1(\as2650.r123[1][6] ),
    .A2(_0815_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4976_ (.A1(_0713_),
    .A2(_0814_),
    .B(_0818_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4977_ (.A1(\as2650.r123[1][7] ),
    .A2(_0815_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4978_ (.A1(_0795_),
    .A2(_0814_),
    .B(_0819_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4979_ (.I(_3551_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4980_ (.A1(_0820_),
    .A2(_3533_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4981_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4982_ (.A1(\as2650.halted ),
    .A2(_3519_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4983_ (.A1(_3483_),
    .A2(_0823_),
    .A3(_3552_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4984_ (.A1(_3484_),
    .A2(_0823_),
    .A3(_3562_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4985_ (.A1(_0800_),
    .A2(_0824_),
    .B(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4986_ (.A1(_0822_),
    .A2(_0826_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4988_ (.I(_0825_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4989_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_3542_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4991_ (.A1(_0831_),
    .A2(_0313_),
    .A3(_0315_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4992_ (.A1(_3483_),
    .A2(_0823_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4993_ (.A1(_3618_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4995_ (.I(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4996_ (.A1(_0832_),
    .A2(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4997_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_0799_),
    .A2(_0835_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4999_ (.I(_0839_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5000_ (.I(_0840_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5001_ (.A1(_3640_),
    .A2(_0824_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5002_ (.A1(_3583_),
    .A2(_0824_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5003_ (.I(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5004_ (.A1(_3572_),
    .A2(_0824_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5005_ (.I(_0845_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5006_ (.A1(_3666_),
    .A2(_0846_),
    .B(_0844_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5007_ (.A1(_3677_),
    .A2(_0835_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5008_ (.A1(_3692_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5009_ (.A1(_3708_),
    .A2(_0844_),
    .B1(_0847_),
    .B2(_0849_),
    .C(_0842_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5010_ (.A1(_3664_),
    .A2(_0842_),
    .B(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5011_ (.A1(_0832_),
    .A2(_0836_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5012_ (.A1(_3715_),
    .A2(_0840_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5013_ (.A1(_0841_),
    .A2(_0851_),
    .B(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5014_ (.A1(_3721_),
    .A2(_0836_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5016_ (.A1(_3731_),
    .A2(_0838_),
    .B(_0854_),
    .C(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5017_ (.I(_0836_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5018_ (.A1(_3721_),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5019_ (.I(_0823_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5020_ (.A1(_3484_),
    .A2(_3537_),
    .A3(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5021_ (.I(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5022_ (.A1(_3740_),
    .A2(_0859_),
    .B(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5023_ (.A1(_0857_),
    .A2(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_3742_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5025_ (.I(_3684_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5026_ (.I(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5027_ (.A1(_3511_),
    .A2(_0833_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5028_ (.I(_0868_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5029_ (.A1(_0865_),
    .A2(_0867_),
    .A3(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5030_ (.I(_0829_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5031_ (.A1(_0864_),
    .A2(_0870_),
    .B(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5032_ (.A1(_3796_),
    .A2(_0830_),
    .B(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5033_ (.I(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5034_ (.I(_0827_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5035_ (.I(_0862_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5037_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_0875_),
    .B(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5038_ (.A1(_0828_),
    .A2(_0874_),
    .B(_0878_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5039_ (.I(_0859_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5040_ (.I(_0840_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5041_ (.I(_0852_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5042_ (.I(_0881_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5043_ (.I(_3852_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5044_ (.A1(_3598_),
    .A2(_0835_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5045_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5046_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5047_ (.I(_3874_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_3855_),
    .A2(_0834_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5049_ (.I(_0888_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5050_ (.I(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5051_ (.I(_0884_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5052_ (.I(_0845_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_0888_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5054_ (.I(_3883_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_0894_),
    .A2(_0846_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5056_ (.A1(_3881_),
    .A2(_0892_),
    .B(_0893_),
    .C(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5057_ (.A1(_0887_),
    .A2(_0890_),
    .B(_0891_),
    .C(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5058_ (.I(_0839_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5059_ (.A1(_0883_),
    .A2(_0886_),
    .B(_0897_),
    .C(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5060_ (.A1(_3843_),
    .A2(_0880_),
    .B(_0882_),
    .C(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5061_ (.A1(_3900_),
    .A2(_0838_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5062_ (.A1(_0879_),
    .A2(_0900_),
    .A3(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5063_ (.I(_0855_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5064_ (.A1(_3908_),
    .A2(_0903_),
    .B(_0869_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5065_ (.I(_3702_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5066_ (.A1(_3842_),
    .A2(_3714_),
    .A3(_0867_),
    .A4(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5067_ (.I(_0861_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5068_ (.I(_3843_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5069_ (.A1(_0908_),
    .A2(_0867_),
    .B1(_0905_),
    .B2(_3742_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5070_ (.A1(_0907_),
    .A2(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5071_ (.A1(_0902_),
    .A2(_0904_),
    .B1(_0906_),
    .B2(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5072_ (.A1(_0830_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5073_ (.A1(_3833_),
    .A2(_0830_),
    .B(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5074_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_0875_),
    .B(_0877_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5075_ (.A1(_0828_),
    .A2(_0913_),
    .B(_0914_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5076_ (.A1(_3835_),
    .A2(_3702_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5077_ (.A1(_3713_),
    .A2(_3868_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5078_ (.A1(_0915_),
    .A2(_0916_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5079_ (.A1(_0279_),
    .A2(_0866_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5080_ (.A1(_0917_),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5081_ (.A1(_0906_),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5082_ (.A1(_0906_),
    .A2(_0919_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5083_ (.A1(_0869_),
    .A2(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5084_ (.A1(_0284_),
    .A2(_0848_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5085_ (.A1(_0288_),
    .A2(_0848_),
    .B(_0889_),
    .C(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5086_ (.A1(_0306_),
    .A2(_0889_),
    .B(_0884_),
    .C(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5087_ (.A1(_3708_),
    .A2(_0885_),
    .B(_0925_),
    .C(_0839_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5088_ (.A1(_0280_),
    .A2(_0898_),
    .B(_0881_),
    .C(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5089_ (.A1(_0321_),
    .A2(_0837_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5090_ (.A1(_0859_),
    .A2(_0927_),
    .A3(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5091_ (.A1(_0277_),
    .A2(_0859_),
    .B(_0862_),
    .C(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5092_ (.A1(_0920_),
    .A2(_0922_),
    .B(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5093_ (.I0(_0266_),
    .I1(_0931_),
    .S(_0829_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5094_ (.I(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5095_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_0875_),
    .B(_0877_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5096_ (.A1(_0828_),
    .A2(_0933_),
    .B(_0934_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(_0822_),
    .A2(_0826_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5098_ (.A1(_0434_),
    .A2(_0346_),
    .B1(_0365_),
    .B2(_0366_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5099_ (.I(_0312_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5100_ (.I(_3548_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5101_ (.I(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5102_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5103_ (.A1(_0937_),
    .A2(_0940_),
    .A3(_3561_),
    .A4(_0833_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5104_ (.I(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5105_ (.I(_0868_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5106_ (.I(\as2650.r123_2[0][3] ),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5107_ (.I(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(_3713_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5109_ (.A1(_3699_),
    .A2(_3867_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5110_ (.A1(_0295_),
    .A2(_3684_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5111_ (.A1(\as2650.r0[2] ),
    .A2(\as2650.r123_2[0][1] ),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5112_ (.A1(_0947_),
    .A2(_0948_),
    .A3(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5113_ (.A1(_0946_),
    .A2(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5114_ (.A1(_0915_),
    .A2(_0916_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5115_ (.A1(_0279_),
    .A2(_0866_),
    .A3(_0917_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5116_ (.A1(_0952_),
    .A2(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5117_ (.A1(_0951_),
    .A2(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5118_ (.A1(_0920_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5119_ (.A1(_0384_),
    .A2(_0848_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5120_ (.A1(_0388_),
    .A2(_0846_),
    .B(_0843_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5121_ (.A1(_0402_),
    .A2(_0844_),
    .B1(_0957_),
    .B2(_0958_),
    .C(_0842_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5122_ (.I(_3930_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5123_ (.A1(_0960_),
    .A2(_0885_),
    .B(_0839_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5124_ (.A1(_0407_),
    .A2(_0840_),
    .B1(_0959_),
    .B2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5125_ (.A1(_0838_),
    .A2(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5126_ (.A1(_0380_),
    .A2(_0838_),
    .B(_0855_),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5127_ (.A1(_0376_),
    .A2(_0856_),
    .B(_0869_),
    .C(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5128_ (.A1(_0943_),
    .A2(_0956_),
    .B(_0965_),
    .C(_0942_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5129_ (.A1(_0936_),
    .A2(_0942_),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5130_ (.A1(_0935_),
    .A2(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5131_ (.I(_0827_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5132_ (.I(_0876_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5133_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_0969_),
    .B(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5134_ (.A1(_0968_),
    .A2(_0971_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5135_ (.I0(_0445_),
    .I1(_0462_),
    .S(_0338_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5136_ (.I(_3604_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5137_ (.I(_3608_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5138_ (.A1(_0973_),
    .A2(_0974_),
    .A3(_0858_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5139_ (.I(_0495_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5140_ (.I(_0845_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_0976_),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5142_ (.A1(_0494_),
    .A2(_0892_),
    .B(_0893_),
    .C(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5143_ (.A1(_0663_),
    .A2(_0890_),
    .B(_0891_),
    .C(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5144_ (.A1(_0307_),
    .A2(_0842_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5145_ (.A1(_0841_),
    .A2(_0980_),
    .A3(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5146_ (.A1(_0492_),
    .A2(_0880_),
    .B(_0975_),
    .C(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5147_ (.A1(_0491_),
    .A2(_0882_),
    .B(_0879_),
    .C(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5148_ (.A1(_0517_),
    .A2(_0903_),
    .B(_0943_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_0920_),
    .A2(_0955_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5150_ (.A1(_0952_),
    .A2(_0953_),
    .B(_0951_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5151_ (.A1(_3712_),
    .A2(_0945_),
    .A3(_0950_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5152_ (.A1(_0947_),
    .A2(_0949_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5153_ (.A1(_0947_),
    .A2(_0949_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5154_ (.A1(_0948_),
    .A2(_0989_),
    .B(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5155_ (.I(\as2650.r123_2[0][4] ),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5156_ (.A1(_3712_),
    .A2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5157_ (.A1(_0991_),
    .A2(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5158_ (.A1(_0991_),
    .A2(_0993_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(_0994_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5160_ (.A1(_3834_),
    .A2(_0944_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(_0390_),
    .A2(\as2650.r123_2[0][0] ),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5162_ (.I(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(\as2650.r0[3] ),
    .A2(\as2650.r123_2[0][2] ),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5164_ (.A1(_0949_),
    .A2(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5165_ (.A1(_0294_),
    .A2(\as2650.r123_2[0][1] ),
    .B1(_3867_),
    .B2(\as2650.r0[2] ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5166_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5167_ (.A1(_0999_),
    .A2(_1003_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5168_ (.A1(_0997_),
    .A2(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5169_ (.A1(_0988_),
    .A2(_0996_),
    .A3(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5170_ (.A1(_0987_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5171_ (.I(_1006_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5172_ (.A1(_0920_),
    .A2(_0955_),
    .A3(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5173_ (.A1(_0868_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5174_ (.A1(_0986_),
    .A2(_1007_),
    .B(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5175_ (.A1(_0984_),
    .A2(_0985_),
    .B(_1011_),
    .C(_0941_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5176_ (.A1(_0972_),
    .A2(_0942_),
    .B(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5177_ (.A1(_0935_),
    .A2(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5178_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_0969_),
    .B(_0970_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5179_ (.A1(_1014_),
    .A2(_1015_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5180_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_0969_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5181_ (.I(_0560_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5182_ (.A1(_0580_),
    .A2(_0977_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5183_ (.A1(_0576_),
    .A2(_0892_),
    .B(_0893_),
    .C(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5184_ (.A1(_0706_),
    .A2(_0890_),
    .B(_0891_),
    .C(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5185_ (.A1(_0561_),
    .A2(_0886_),
    .B(_1020_),
    .C(_0898_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5186_ (.A1(_1017_),
    .A2(_0880_),
    .B(_0882_),
    .C(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5187_ (.I(_3847_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5188_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5189_ (.I(_3849_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5190_ (.A1(_1024_),
    .A2(_1025_),
    .A3(_0588_),
    .A4(_0858_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5191_ (.A1(_1022_),
    .A2(_1026_),
    .B(_0903_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5192_ (.A1(_0559_),
    .A2(_0903_),
    .B(_0943_),
    .C(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5193_ (.A1(_0987_),
    .A2(_1008_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5194_ (.A1(_0988_),
    .A2(_1005_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5195_ (.A1(_0988_),
    .A2(_1005_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5196_ (.A1(_0996_),
    .A2(_1030_),
    .B(_1031_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5197_ (.A1(_3699_),
    .A2(_0944_),
    .A3(_1004_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5198_ (.A1(_3859_),
    .A2(\as2650.r123_2[0][3] ),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5199_ (.A1(\as2650.r0[5] ),
    .A2(\as2650.r123_2[0][0] ),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5200_ (.A1(\as2650.r0[4] ),
    .A2(\as2650.r123_2[0][1] ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5201_ (.A1(_1000_),
    .A2(_1035_),
    .A3(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5202_ (.A1(_1034_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5203_ (.I(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5204_ (.A1(_1033_),
    .A2(_1039_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5205_ (.A1(_0999_),
    .A2(_1003_),
    .B(_1001_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_3681_),
    .A2(\as2650.r123_2[0][5] ),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5207_ (.A1(_1041_),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5208_ (.A1(_3834_),
    .A2(\as2650.r123_2[0][4] ),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5209_ (.A1(_1043_),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5210_ (.A1(_1040_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5211_ (.A1(_1032_),
    .A2(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5212_ (.A1(_0994_),
    .A2(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5213_ (.A1(_1029_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5214_ (.A1(_1009_),
    .A2(_1049_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5215_ (.A1(_0876_),
    .A2(_1050_),
    .B(_0871_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5216_ (.A1(_0553_),
    .A2(_0942_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5217_ (.A1(_1028_),
    .A2(_1051_),
    .B(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5218_ (.A1(_0935_),
    .A2(_1053_),
    .B(_0970_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5219_ (.A1(_1016_),
    .A2(_1054_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5220_ (.I(_0711_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5221_ (.A1(_1029_),
    .A2(_1048_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5222_ (.A1(_1009_),
    .A2(_1049_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5223_ (.A1(_1056_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5224_ (.A1(_1041_),
    .A2(_1042_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5225_ (.A1(_1043_),
    .A2(_1044_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5226_ (.A1(_1059_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5227_ (.I(_1040_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5228_ (.A1(_1033_),
    .A2(_1039_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5229_ (.A1(_1062_),
    .A2(_1045_),
    .B(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5230_ (.A1(_1034_),
    .A2(_1037_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5231_ (.A1(_3711_),
    .A2(\as2650.r123_2[0][6] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(_0296_),
    .A2(_0944_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5233_ (.A1(_0498_),
    .A2(_3702_),
    .B1(_3868_),
    .B2(_0390_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5234_ (.I(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5235_ (.A1(_0498_),
    .A2(_3867_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5236_ (.A1(_1036_),
    .A2(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(_1069_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(\as2650.r0[6] ),
    .A2(_3684_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5239_ (.A1(_1072_),
    .A2(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5240_ (.A1(_1066_),
    .A2(_1067_),
    .A3(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5241_ (.A1(_1065_),
    .A2(_1075_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5242_ (.I(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5243_ (.I(_1035_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(_1000_),
    .A2(_1036_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5245_ (.A1(_1000_),
    .A2(_1036_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5246_ (.A1(_1078_),
    .A2(_1079_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5247_ (.A1(_3835_),
    .A2(_0501_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5248_ (.A1(_1081_),
    .A2(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(_1081_),
    .A2(_1082_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5250_ (.A1(_1083_),
    .A2(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5251_ (.A1(_0278_),
    .A2(_0992_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5252_ (.A1(_1085_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5253_ (.A1(_1077_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5254_ (.A1(_1061_),
    .A2(_1064_),
    .A3(_1088_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5255_ (.A1(_0994_),
    .A2(_1047_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5256_ (.A1(_1032_),
    .A2(_1046_),
    .B(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5257_ (.A1(_1089_),
    .A2(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_1089_),
    .A2(_1091_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5259_ (.A1(_1092_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5260_ (.A1(_1058_),
    .A2(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5261_ (.I(_0507_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5262_ (.I(_0669_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5263_ (.I(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5264_ (.A1(_0667_),
    .A2(_0977_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5265_ (.A1(_1098_),
    .A2(_0892_),
    .B(_0844_),
    .C(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5266_ (.I(_0720_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5267_ (.A1(_1101_),
    .A2(_0890_),
    .B(_0891_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5268_ (.A1(_1096_),
    .A2(_0886_),
    .B1(_1100_),
    .B2(_1102_),
    .C(_0898_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5269_ (.A1(_0662_),
    .A2(_0880_),
    .B(_0881_),
    .C(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5270_ (.A1(_1024_),
    .A2(_1025_),
    .A3(_0679_),
    .A4(_0858_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5271_ (.A1(_1104_),
    .A2(_1105_),
    .B(_0856_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5272_ (.A1(_0660_),
    .A2(_0856_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5273_ (.A1(_0907_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5274_ (.A1(_0876_),
    .A2(_1095_),
    .B1(_1106_),
    .B2(_1108_),
    .C(_0871_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5275_ (.A1(_1055_),
    .A2(_0830_),
    .B(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5276_ (.A1(_0935_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5277_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_0969_),
    .B(_0970_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5278_ (.A1(_1111_),
    .A2(_1112_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5279_ (.I(_3645_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5280_ (.I(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5281_ (.I(_0781_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1115_),
    .A2(_0846_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5283_ (.A1(_0780_),
    .A2(_0977_),
    .B(_0889_),
    .C(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5284_ (.A1(_0776_),
    .A2(_0893_),
    .B(_0885_),
    .C(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5285_ (.A1(_0775_),
    .A2(_0886_),
    .B(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5286_ (.A1(_0841_),
    .A2(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5287_ (.A1(_1114_),
    .A2(_0841_),
    .B(_0881_),
    .C(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5288_ (.A1(_0790_),
    .A2(_0882_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5289_ (.A1(_0774_),
    .A2(_0879_),
    .B(_0862_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5290_ (.A1(_0879_),
    .A2(_1122_),
    .B(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5291_ (.A1(_1058_),
    .A2(_1094_),
    .B(_1092_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5292_ (.A1(_1065_),
    .A2(_1075_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5293_ (.A1(_1077_),
    .A2(_1087_),
    .B(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5294_ (.A1(_0392_),
    .A2(_0945_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5295_ (.A1(_3836_),
    .A2(\as2650.r123_2[0][6] ),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5296_ (.A1(_1128_),
    .A2(_1129_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5297_ (.A1(_1085_),
    .A2(_1086_),
    .B(_1083_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5298_ (.A1(_1066_),
    .A2(_1067_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_1066_),
    .A2(_1067_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5300_ (.A1(_1132_),
    .A2(_1133_),
    .A3(_1074_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5301_ (.A1(_1068_),
    .A2(_1073_),
    .B(_1071_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5302_ (.A1(_3713_),
    .A2(\as2650.r123_2[0][7] ),
    .A3(_1132_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5303_ (.A1(\as2650.r123_2[0][7] ),
    .A2(_1132_),
    .B(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5304_ (.A1(\as2650.r0[7] ),
    .A2(_0866_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5305_ (.A1(_0278_),
    .A2(_0501_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5306_ (.A1(_1070_),
    .A2(_1138_),
    .A3(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5307_ (.A1(_1137_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5308_ (.A1(_1134_),
    .A2(_1135_),
    .A3(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5309_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5310_ (.A1(_1127_),
    .A2(_1143_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5311_ (.A1(_1064_),
    .A2(_1088_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5312_ (.A1(_1064_),
    .A2(_1088_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5313_ (.A1(_1061_),
    .A2(_1145_),
    .B(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5314_ (.A1(_0406_),
    .A2(_0992_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5315_ (.A1(_0661_),
    .A2(_0905_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5316_ (.A1(_1147_),
    .A2(_1148_),
    .A3(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5317_ (.A1(_1125_),
    .A2(_1144_),
    .A3(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5318_ (.A1(_0907_),
    .A2(_1151_),
    .B(_0829_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5319_ (.A1(_1124_),
    .A2(_1152_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5320_ (.I(_0741_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5321_ (.A1(_1154_),
    .A2(_0871_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5322_ (.A1(_1153_),
    .A2(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_0875_),
    .B(_0877_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5324_ (.A1(_0828_),
    .A2(_1156_),
    .B(_1157_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5325_ (.I(_0803_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5326_ (.I(_3534_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5327_ (.A1(_1158_),
    .A2(_1159_),
    .A3(_0826_),
    .A4(_0907_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5328_ (.I(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5329_ (.I(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5330_ (.A1(_0867_),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5331_ (.A1(_0874_),
    .A2(_1162_),
    .B(_1163_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5332_ (.I(_1160_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(_0905_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5334_ (.A1(_0913_),
    .A2(_1162_),
    .B(_1165_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5335_ (.A1(_3868_),
    .A2(_1164_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5336_ (.A1(_0933_),
    .A2(_1162_),
    .B(_1166_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5337_ (.I0(_0967_),
    .I1(_0945_),
    .S(_1164_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5338_ (.I(_1167_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5339_ (.I0(_1013_),
    .I1(_0992_),
    .S(_1164_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5340_ (.I(_1168_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5341_ (.I0(_1053_),
    .I1(_0501_),
    .S(_1161_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_1169_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5343_ (.I0(_1110_),
    .I1(\as2650.r123_2[0][6] ),
    .S(_1161_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5344_ (.I(_1170_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5345_ (.A1(_1153_),
    .A2(_1155_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5346_ (.I0(_1171_),
    .I1(\as2650.r123_2[0][7] ),
    .S(_1161_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5347_ (.I(_1172_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5348_ (.I(\as2650.r123[3][0] ),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5349_ (.I(_1173_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5350_ (.I(\as2650.r123[3][1] ),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5351_ (.I(_1174_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5352_ (.I(\as2650.r123[3][2] ),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_1175_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5354_ (.I(\as2650.r123[3][3] ),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5355_ (.I(_1176_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5356_ (.I(\as2650.r123[3][4] ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5357_ (.I(_1177_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5358_ (.I(\as2650.r123[3][5] ),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5359_ (.I(_1178_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(\as2650.r123[3][6] ),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5361_ (.I(_1179_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(\as2650.r123[3][7] ),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5363_ (.I(_1180_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5364_ (.A1(_0820_),
    .A2(_0826_),
    .B(_0943_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5365_ (.I(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5366_ (.I(_1181_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5367_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_1183_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5368_ (.A1(_0874_),
    .A2(_1182_),
    .B(_1184_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5369_ (.A1(\as2650.r123_2[1][1] ),
    .A2(_1183_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5370_ (.A1(_0913_),
    .A2(_1182_),
    .B(_1185_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5371_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_1183_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5372_ (.A1(_0933_),
    .A2(_1182_),
    .B(_1186_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5373_ (.I(_1181_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5374_ (.I0(_0967_),
    .I1(\as2650.r123_2[1][3] ),
    .S(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5375_ (.I(_1188_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5376_ (.I0(_1013_),
    .I1(\as2650.r123_2[1][4] ),
    .S(_1187_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_1189_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5378_ (.I0(_1053_),
    .I1(\as2650.r123_2[1][5] ),
    .S(_1187_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5379_ (.I(_1190_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5380_ (.I0(_1110_),
    .I1(\as2650.r123_2[1][6] ),
    .S(_1187_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5381_ (.I(_1191_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_1183_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5383_ (.A1(_1156_),
    .A2(_1182_),
    .B(_1192_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5384_ (.I(\as2650.psu[5] ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5385_ (.I(_3530_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5386_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5387_ (.A1(_0820_),
    .A2(_3497_),
    .A3(_3535_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5388_ (.I(_3575_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5389_ (.A1(_3496_),
    .A2(_3504_),
    .A3(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5390_ (.I(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5391_ (.A1(_3536_),
    .A2(_1196_),
    .A3(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5392_ (.I(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5393_ (.A1(_1195_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_3576_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5395_ (.I(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5396_ (.I(_3573_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5397_ (.I(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5398_ (.A1(_1206_),
    .A2(_3674_),
    .A3(_3935_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5399_ (.I(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_3565_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_1209_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5402_ (.I(_1210_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5403_ (.A1(_0822_),
    .A2(_1208_),
    .B(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(_1204_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5405_ (.I(_0547_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5406_ (.A1(_1205_),
    .A2(_1197_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5410_ (.I(\as2650.psl[7] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5411_ (.A1(_1219_),
    .A2(_3496_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5412_ (.A1(\as2650.psl[6] ),
    .A2(_0820_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5413_ (.A1(_1220_),
    .A2(_1221_),
    .B(_0822_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5414_ (.A1(_1195_),
    .A2(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5415_ (.A1(_1214_),
    .A2(_1218_),
    .A3(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5416_ (.A1(_1202_),
    .A2(_1213_),
    .B(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5417_ (.A1(_1194_),
    .A2(_1199_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5418_ (.A1(_1158_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5419_ (.I(_0802_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5420_ (.I(_1198_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5421_ (.A1(_1228_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5422_ (.I(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5423_ (.A1(_3490_),
    .A2(_1209_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5425_ (.I(_3593_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5426_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(_1235_),
    .A2(_3848_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5429_ (.A1(_3528_),
    .A2(_3544_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5430_ (.I(_1238_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5431_ (.A1(_3671_),
    .A2(_1239_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5432_ (.I(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5433_ (.A1(_1237_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5434_ (.I(_1242_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5435_ (.I(_3573_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5436_ (.A1(_3752_),
    .A2(_3499_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5437_ (.A1(_1244_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5438_ (.A1(_1246_),
    .A2(_3581_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5439_ (.I(\as2650.halted ),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5440_ (.A1(_3527_),
    .A2(_3589_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_1249_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5442_ (.A1(_3672_),
    .A2(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5443_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5444_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5445_ (.A1(_1248_),
    .A2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5446_ (.I(_1211_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5447_ (.I(_1207_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5448_ (.A1(_1228_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5449_ (.A1(_3497_),
    .A2(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5450_ (.A1(_1255_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5451_ (.A1(_1243_),
    .A2(_1247_),
    .A3(_1254_),
    .A4(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5452_ (.A1(_3510_),
    .A2(_1231_),
    .A3(_1233_),
    .A4(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5453_ (.A1(_1225_),
    .A2(_1227_),
    .A3(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5454_ (.I(_1203_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5455_ (.I(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5456_ (.I(_3490_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5457_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5458_ (.I(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5459_ (.A1(_1017_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5460_ (.I(_0579_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5461_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5462_ (.I(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5463_ (.I(_1195_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5464_ (.I(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5465_ (.A1(_3553_),
    .A2(_1208_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5466_ (.A1(_1270_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5467_ (.A1(\as2650.psu[5] ),
    .A2(_1271_),
    .B(_1273_),
    .C(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5468_ (.A1(_1268_),
    .A2(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5469_ (.A1(_1264_),
    .A2(_1277_),
    .B(_1262_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_3519_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5472_ (.A1(_1193_),
    .A2(_1262_),
    .B(_1278_),
    .C(_1280_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5473_ (.A1(_0737_),
    .A2(_0727_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5474_ (.A1(_0727_),
    .A2(_3661_),
    .B(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5475_ (.A1(_0261_),
    .A2(_0353_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5476_ (.I(_3805_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5477_ (.A1(_1284_),
    .A2(_3813_),
    .B1(_3818_),
    .B2(_3761_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5478_ (.A1(_3921_),
    .A2(_0346_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5479_ (.A1(_0344_),
    .A2(_1283_),
    .B1(_1285_),
    .B2(_1286_),
    .C(_0446_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(_0445_),
    .A2(_0534_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5481_ (.I(_0695_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5482_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_1287_),
    .B2(_1288_),
    .C(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5483_ (.A1(_0692_),
    .A2(_0731_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5484_ (.I(\as2650.psl[1] ),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5485_ (.A1(_0705_),
    .A2(_0718_),
    .A3(_0723_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5486_ (.A1(_1292_),
    .A2(_0718_),
    .B(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5487_ (.A1(_0736_),
    .A2(_1282_),
    .B1(_1290_),
    .B2(_1291_),
    .C(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5488_ (.A1(_0736_),
    .A2(_1282_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5489_ (.A1(_1292_),
    .A2(_0718_),
    .A3(_1296_),
    .B(_0572_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5490_ (.A1(_1295_),
    .A2(_1297_),
    .B(_1273_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5491_ (.I(_1267_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5492_ (.A1(_1299_),
    .A2(_3818_),
    .A3(_1288_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5493_ (.A1(_3764_),
    .A2(_1286_),
    .A3(_1291_),
    .A4(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5494_ (.A1(_1298_),
    .A2(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5495_ (.A1(_3833_),
    .A2(_0266_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5496_ (.A1(_3796_),
    .A2(_0936_),
    .A3(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5497_ (.A1(_0465_),
    .A2(_0553_),
    .A3(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5498_ (.A1(_1055_),
    .A2(_1305_),
    .B(_1154_),
    .C(_0572_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5499_ (.I(_1299_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5500_ (.I(_3566_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5501_ (.I(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5502_ (.A1(_3934_),
    .A2(_1309_),
    .A3(_3574_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5503_ (.I(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5504_ (.A1(_1101_),
    .A2(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5505_ (.A1(_0280_),
    .A2(_3842_),
    .A3(_3715_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5506_ (.A1(_0662_),
    .A2(_0560_),
    .A3(_0492_),
    .A4(_0407_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5507_ (.A1(_1313_),
    .A2(_1314_),
    .B(_1113_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5508_ (.A1(_0769_),
    .A2(_1312_),
    .B1(_1315_),
    .B2(_1311_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5509_ (.A1(_1307_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5510_ (.I(_1308_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5511_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5512_ (.I(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5513_ (.A1(_1302_),
    .A2(_1306_),
    .B(_1317_),
    .C(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5514_ (.I(_1255_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5515_ (.I(_3530_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5516_ (.I(_1323_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5517_ (.A1(_3611_),
    .A2(_1215_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5518_ (.I(_1325_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5519_ (.A1(_0312_),
    .A2(_1324_),
    .A3(_1247_),
    .A4(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(_1309_),
    .A2(_1323_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5521_ (.A1(_3673_),
    .A2(_3548_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5522_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5523_ (.I(_0311_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5524_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5525_ (.A1(_3628_),
    .A2(_1310_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5526_ (.A1(_3541_),
    .A2(_0358_),
    .A3(_3552_),
    .A4(_3810_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5527_ (.A1(_3529_),
    .A2(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5528_ (.A1(_1333_),
    .A2(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5529_ (.A1(_1332_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5530_ (.I(_3512_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5531_ (.A1(_3593_),
    .A2(_3499_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5532_ (.I(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5533_ (.A1(_3671_),
    .A2(_1239_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5534_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5535_ (.A1(_1338_),
    .A2(_1263_),
    .A3(_1340_),
    .A4(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5536_ (.A1(_1203_),
    .A2(_1247_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5537_ (.A1(_1214_),
    .A2(_1237_),
    .A3(_1212_),
    .A4(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5538_ (.A1(_1330_),
    .A2(_1337_),
    .A3(_1343_),
    .A4(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5539_ (.A1(_1322_),
    .A2(_1327_),
    .B(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5540_ (.A1(_3509_),
    .A2(_1199_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5541_ (.A1(_1203_),
    .A2(_1247_),
    .A3(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5542_ (.A1(_1196_),
    .A2(_1349_),
    .B(_3577_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5543_ (.I(_3673_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5544_ (.I(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5545_ (.A1(_1228_),
    .A2(_1352_),
    .A3(_1207_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5546_ (.A1(_3537_),
    .A2(_1350_),
    .A3(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5547_ (.A1(_3569_),
    .A2(_3934_),
    .A3(_3585_),
    .A4(_3787_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5548_ (.A1(_1235_),
    .A2(_1323_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5549_ (.A1(_1355_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5550_ (.A1(_3529_),
    .A2(_3673_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(_1308_),
    .A2(_1209_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5552_ (.I(_1359_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5553_ (.A1(_3672_),
    .A2(_1250_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5554_ (.I(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5555_ (.A1(_3676_),
    .A2(_1358_),
    .B(_1360_),
    .C(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5556_ (.A1(_1309_),
    .A2(_1265_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5557_ (.I(_3618_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5558_ (.A1(_1365_),
    .A2(_0799_),
    .B1(_1334_),
    .B2(_3490_),
    .C(\as2650.halted ),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5559_ (.A1(_0359_),
    .A2(_1245_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5560_ (.A1(_3595_),
    .A2(_3491_),
    .B(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5561_ (.A1(_0727_),
    .A2(_1364_),
    .B(_1366_),
    .C(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5562_ (.A1(_1357_),
    .A2(_1363_),
    .A3(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5563_ (.A1(_1354_),
    .A2(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5564_ (.A1(_1347_),
    .A2(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5565_ (.I(_0937_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5566_ (.I(_1373_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5567_ (.A1(_0707_),
    .A2(_1246_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5568_ (.I(_3595_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_1355_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5570_ (.A1(_1376_),
    .A2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5571_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5572_ (.I(_0661_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5573_ (.A1(_1380_),
    .A2(_1229_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5574_ (.I(_3491_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5575_ (.I(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5576_ (.A1(_1229_),
    .A2(_1315_),
    .B(_1381_),
    .C(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(_1194_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5578_ (.I(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_1098_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5580_ (.I(\as2650.psl[6] ),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5581_ (.A1(_1388_),
    .A2(_1387_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5582_ (.A1(_3534_),
    .A2(_1387_),
    .B(_1257_),
    .C(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5583_ (.A1(_0707_),
    .A2(_1377_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5584_ (.I(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5585_ (.A1(_1386_),
    .A2(_1390_),
    .B(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5586_ (.A1(_3597_),
    .A2(_0775_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5587_ (.I(_3597_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5588_ (.A1(_1395_),
    .A2(_3664_),
    .A3(_0656_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5589_ (.A1(_1384_),
    .A2(_1393_),
    .B(_1394_),
    .C(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5590_ (.I(_1378_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5591_ (.A1(_1398_),
    .A2(_0776_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_1378_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5593_ (.I(_3661_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5594_ (.A1(_3816_),
    .A2(_0887_),
    .A3(_0307_),
    .A4(_0449_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5595_ (.A1(_1400_),
    .A2(_1401_),
    .A3(_1402_),
    .A4(_0768_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5596_ (.A1(_1379_),
    .A2(_1397_),
    .B(_1399_),
    .C(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5597_ (.A1(_1375_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5598_ (.I(_0781_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5599_ (.I(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5600_ (.I(_1407_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5601_ (.I(_3675_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5602_ (.I(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_1408_),
    .A2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5604_ (.I(_3666_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5605_ (.I(_1412_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5606_ (.I(_1413_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5607_ (.I(_0894_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5608_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5609_ (.I(_0286_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5610_ (.I(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5611_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5612_ (.I(_0388_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5613_ (.I(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5614_ (.A1(_1414_),
    .A2(_1416_),
    .A3(_1419_),
    .A4(_1421_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5615_ (.I(_0976_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5616_ (.I(_1387_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5618_ (.A1(_1423_),
    .A2(_1271_),
    .A3(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5619_ (.A1(_1410_),
    .A2(_1422_),
    .A3(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5620_ (.A1(_1374_),
    .A2(_1405_),
    .A3(_1411_),
    .A4(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5621_ (.A1(_1372_),
    .A2(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5622_ (.I(_3513_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5623_ (.I(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5624_ (.A1(_1388_),
    .A2(_1372_),
    .B(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5625_ (.A1(_1321_),
    .A2(_1429_),
    .B(_1432_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5626_ (.I(_1332_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5627_ (.I(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5628_ (.A1(_3829_),
    .A2(_0730_),
    .A3(_0734_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5629_ (.A1(_0338_),
    .A2(_0731_),
    .B1(_1435_),
    .B2(_0739_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5630_ (.A1(_3560_),
    .A2(_1436_),
    .B(_1298_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5631_ (.I(_1324_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5632_ (.I(_1438_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5633_ (.I(_1439_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5634_ (.A1(_1114_),
    .A2(_1311_),
    .B(_1312_),
    .C(_1440_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5635_ (.I(_1373_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5636_ (.A1(_1442_),
    .A2(_1411_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_1377_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5638_ (.I(_1444_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5639_ (.I(_1267_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5640_ (.A1(_1113_),
    .A2(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5641_ (.I(_1406_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5642_ (.I(_1448_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5643_ (.A1(\as2650.psl[7] ),
    .A2(_1407_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5644_ (.A1(_1159_),
    .A2(_1449_),
    .B(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5645_ (.A1(_0802_),
    .A2(_1206_),
    .A3(_3674_),
    .A4(_3815_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5646_ (.I(_3667_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5647_ (.I(net2),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5648_ (.I(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5649_ (.I(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5650_ (.I(\as2650.psl[5] ),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5651_ (.I(_3882_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5652_ (.I(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5653_ (.I(_1459_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5654_ (.A1(_1219_),
    .A2(_0782_),
    .B1(_0495_),
    .B2(_3650_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5655_ (.A1(\as2650.psl[1] ),
    .A2(_1460_),
    .B1(_0288_),
    .B2(\as2650.overflow ),
    .C(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5656_ (.A1(_3644_),
    .A2(_1420_),
    .B1(_0580_),
    .B2(_1457_),
    .C(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5657_ (.A1(_3767_),
    .A2(_1453_),
    .B1(_1456_),
    .B2(_1388_),
    .C(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5658_ (.A1(_1244_),
    .A2(_1234_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5659_ (.A1(_3542_),
    .A2(_3814_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5660_ (.A1(_1228_),
    .A2(_1465_),
    .A3(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5661_ (.I(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5662_ (.A1(_1406_),
    .A2(_3661_),
    .B1(_0960_),
    .B2(_0286_),
    .C1(_0699_),
    .C2(_1098_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5663_ (.A1(_3667_),
    .A2(_3852_),
    .B1(_0402_),
    .B2(_0976_),
    .C1(_1096_),
    .C2(_1269_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5664_ (.I(net8),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5665_ (.I(_1471_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5666_ (.A1(_1472_),
    .A2(_0306_),
    .B(_1452_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5667_ (.A1(_0894_),
    .A2(_3707_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5668_ (.A1(_1469_),
    .A2(_1470_),
    .A3(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5669_ (.A1(_1452_),
    .A2(_1464_),
    .B(_1468_),
    .C(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5670_ (.I(net9),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(_1477_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5672_ (.I(_1478_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5674_ (.I(\as2650.psu[7] ),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5675_ (.I(\as2650.psu[2] ),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5676_ (.I(net1),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5677_ (.I(\as2650.psu[1] ),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5678_ (.I(net27),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5679_ (.A1(_1484_),
    .A2(_3883_),
    .B1(_0670_),
    .B2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5680_ (.A1(\as2650.psu[3] ),
    .A2(_1472_),
    .B1(_1483_),
    .B2(\as2650.psu[5] ),
    .C(_1486_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5681_ (.A1(_1481_),
    .A2(_1406_),
    .B1(_0286_),
    .B2(_1482_),
    .C(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5682_ (.A1(\as2650.psu[0] ),
    .A2(_1453_),
    .B1(_1480_),
    .B2(\as2650.psu[4] ),
    .C(_1488_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5683_ (.A1(_1467_),
    .A2(_1489_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5684_ (.A1(_1257_),
    .A2(_1476_),
    .A3(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5685_ (.A1(_1257_),
    .A2(_1451_),
    .B(_1491_),
    .C(_1439_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5686_ (.A1(_1447_),
    .A2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5687_ (.A1(_1445_),
    .A2(_1493_),
    .B(_1394_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5688_ (.A1(_1399_),
    .A2(_1494_),
    .B(_1410_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5689_ (.A1(_1434_),
    .A2(_1437_),
    .A3(_1441_),
    .B1(_1443_),
    .B2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5690_ (.A1(\as2650.psl[7] ),
    .A2(_1372_),
    .B(_1431_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5691_ (.A1(_1372_),
    .A2(_1496_),
    .B(_1497_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5692_ (.A1(_1234_),
    .A2(_3566_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5693_ (.A1(_3779_),
    .A2(_1498_),
    .A3(_0821_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5694_ (.A1(_1205_),
    .A2(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5695_ (.A1(_1251_),
    .A2(_1358_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5696_ (.A1(_1500_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5697_ (.I(_3515_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5698_ (.I(_1500_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5699_ (.I(_1504_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5700_ (.A1(_1253_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5701_ (.I(_1351_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5702_ (.A1(_1448_),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5703_ (.A1(_1383_),
    .A2(_1503_),
    .A3(_1506_),
    .A4(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5704_ (.A1(_1502_),
    .A2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5705_ (.I(_1510_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5706_ (.I(_1253_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5707_ (.A1(_1340_),
    .A2(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5708_ (.A1(_1414_),
    .A2(_1512_),
    .B(_1513_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5709_ (.I(_1510_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5710_ (.A1(_1158_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5711_ (.A1(_1511_),
    .A2(_1514_),
    .B(_1516_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5712_ (.A1(_1416_),
    .A2(_1512_),
    .B(_1513_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5713_ (.A1(_3497_),
    .A2(_1515_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5714_ (.A1(_1511_),
    .A2(_1517_),
    .B(_1518_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_1206_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5716_ (.I(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5717_ (.I(_1520_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5718_ (.I(_1362_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5719_ (.A1(_1522_),
    .A2(_1515_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5720_ (.A1(_1521_),
    .A2(_1511_),
    .B1(_1523_),
    .B2(_1419_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5721_ (.I(_1524_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5722_ (.I(_1408_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5723_ (.I(_1507_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5724_ (.I(_1526_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5725_ (.I(_1386_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5727_ (.A1(_1525_),
    .A2(_1527_),
    .B(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5728_ (.A1(_1503_),
    .A2(_1522_),
    .A3(_1530_),
    .B(_1214_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5729_ (.A1(_1271_),
    .A2(_1523_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5730_ (.A1(_1531_),
    .A2(_1532_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5731_ (.A1(_3787_),
    .A2(_1511_),
    .B1(_1523_),
    .B2(_1425_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5732_ (.I(_1533_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5733_ (.A1(_1376_),
    .A2(_1515_),
    .B1(_1523_),
    .B2(_1525_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5734_ (.I(_1534_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5735_ (.I(\as2650.pc[0] ),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5736_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_1536_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5738_ (.I(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5739_ (.I(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5740_ (.I(\as2650.stack_ptr[2] ),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5741_ (.I(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5742_ (.I(\as2650.stack_ptr[1] ),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5743_ (.I(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5744_ (.I(\as2650.stack_ptr[0] ),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5745_ (.A1(_1543_),
    .A2(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_1546_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5748_ (.A1(_3545_),
    .A2(_3547_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5749_ (.I(_1548_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5750_ (.A1(_1205_),
    .A2(_3594_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5751_ (.A1(_3524_),
    .A2(_1466_),
    .A3(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5752_ (.A1(_3594_),
    .A2(_1499_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(_1550_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5754_ (.A1(_1244_),
    .A2(_1351_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5755_ (.I(\as2650.cycle[3] ),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5756_ (.I(\as2650.cycle[2] ),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5757_ (.A1(_1555_),
    .A2(_1556_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5758_ (.A1(_1249_),
    .A2(_1557_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5759_ (.A1(_3600_),
    .A2(_0938_),
    .B1(_1558_),
    .B2(_1551_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5760_ (.A1(_3585_),
    .A2(_3626_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5761_ (.A1(_1554_),
    .A2(_1559_),
    .B(_1560_),
    .C(_0547_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5762_ (.I(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5763_ (.A1(_1549_),
    .A2(_1551_),
    .B1(_1553_),
    .B2(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5764_ (.A1(_3515_),
    .A2(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5765_ (.A1(_1541_),
    .A2(_1547_),
    .A3(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5766_ (.I(_1565_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5768_ (.I(_1566_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5769_ (.A1(\as2650.stack[2][0] ),
    .A2(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5770_ (.A1(_1539_),
    .A2(_1567_),
    .B(_1569_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5771_ (.I(\as2650.pc[1] ),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5772_ (.I(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5773_ (.I(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5774_ (.I(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5775_ (.I(_1565_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5776_ (.I0(_1573_),
    .I1(\as2650.stack[2][1] ),
    .S(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5777_ (.I(_1575_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5778_ (.I(\as2650.pc[2] ),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5779_ (.I(_1576_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5781_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5782_ (.I0(_1579_),
    .I1(\as2650.stack[2][2] ),
    .S(_1574_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5783_ (.I(_1580_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5784_ (.I(\as2650.pc[3] ),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5785_ (.I(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5786_ (.I(_1582_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5787_ (.I(_1566_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(\as2650.stack[2][3] ),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5789_ (.A1(_1583_),
    .A2(_1567_),
    .B(_1585_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5790_ (.I(\as2650.pc[4] ),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5791_ (.I(_1586_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5792_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5794_ (.I(_1566_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5795_ (.I0(_1589_),
    .I1(\as2650.stack[2][4] ),
    .S(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5796_ (.I(_1591_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5797_ (.I(\as2650.pc[5] ),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5798_ (.I(_1592_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5799_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5800_ (.I(_1594_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5801_ (.A1(\as2650.stack[2][5] ),
    .A2(_1584_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5802_ (.A1(_1595_),
    .A2(_1567_),
    .B(_1596_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(\as2650.pc[6] ),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5804_ (.I(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5805_ (.I(_1598_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5806_ (.I(_1599_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(\as2650.stack[2][6] ),
    .A2(_1584_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5808_ (.A1(_1600_),
    .A2(_1567_),
    .B(_1601_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5809_ (.I(\as2650.pc[7] ),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5810_ (.I(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5811_ (.I(_1603_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5812_ (.A1(\as2650.stack[2][7] ),
    .A2(_1584_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5813_ (.A1(_1604_),
    .A2(_1568_),
    .B(_1605_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5814_ (.I(\as2650.pc[8] ),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5815_ (.I(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5816_ (.I(_1607_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5817_ (.I(_1608_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5818_ (.I(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5819_ (.I0(_1610_),
    .I1(\as2650.stack[2][8] ),
    .S(_1590_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5820_ (.I(_1611_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5821_ (.I(\as2650.pc[9] ),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5822_ (.I(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5823_ (.I(_1613_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5824_ (.A1(\as2650.stack[2][9] ),
    .A2(_1574_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5825_ (.A1(_1614_),
    .A2(_1568_),
    .B(_1615_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5826_ (.I(\as2650.pc[10] ),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5827_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(\as2650.stack[2][10] ),
    .A2(_1574_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5829_ (.A1(_1617_),
    .A2(_1568_),
    .B(_1618_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5830_ (.I(\as2650.pc[11] ),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5831_ (.I(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5832_ (.I(_1620_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5833_ (.I(_1621_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5834_ (.I0(_1622_),
    .I1(\as2650.stack[2][11] ),
    .S(_1590_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5835_ (.I(_1623_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5836_ (.I(\as2650.pc[12] ),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5837_ (.I(_1624_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5838_ (.I(_1625_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5839_ (.I0(_1626_),
    .I1(\as2650.stack[2][12] ),
    .S(_1590_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5840_ (.I(_1627_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5841_ (.A1(_1541_),
    .A2(_3515_),
    .A3(_1563_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(_1547_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5843_ (.I(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_1630_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5845_ (.I(_1630_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(\as2650.stack[6][0] ),
    .A2(_1632_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5847_ (.A1(_1539_),
    .A2(_1631_),
    .B(_1633_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5848_ (.I(_1629_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5849_ (.I0(_1573_),
    .I1(\as2650.stack[6][1] ),
    .S(_1634_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5850_ (.I(_1635_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5851_ (.I0(_1579_),
    .I1(\as2650.stack[6][2] ),
    .S(_1634_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5852_ (.I(_1636_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5853_ (.I(_1630_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5854_ (.A1(\as2650.stack[6][3] ),
    .A2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5855_ (.A1(_1583_),
    .A2(_1631_),
    .B(_1638_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5856_ (.I(_1630_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5857_ (.I0(_1589_),
    .I1(\as2650.stack[6][4] ),
    .S(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5858_ (.I(_1640_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5859_ (.A1(\as2650.stack[6][5] ),
    .A2(_1637_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5860_ (.A1(_1595_),
    .A2(_1631_),
    .B(_1641_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5861_ (.A1(\as2650.stack[6][6] ),
    .A2(_1637_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5862_ (.A1(_1600_),
    .A2(_1631_),
    .B(_1642_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5863_ (.A1(\as2650.stack[6][7] ),
    .A2(_1637_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5864_ (.A1(_1604_),
    .A2(_1632_),
    .B(_1643_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5865_ (.I0(_1610_),
    .I1(\as2650.stack[6][8] ),
    .S(_1639_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_1644_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5867_ (.A1(\as2650.stack[6][9] ),
    .A2(_1634_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5868_ (.A1(_1614_),
    .A2(_1632_),
    .B(_1645_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5869_ (.A1(\as2650.stack[6][10] ),
    .A2(_1634_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5870_ (.A1(_1617_),
    .A2(_1632_),
    .B(_1646_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5871_ (.I0(_1622_),
    .I1(\as2650.stack[6][11] ),
    .S(_1639_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5872_ (.I(_1647_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5873_ (.I0(_1626_),
    .I1(\as2650.stack[6][12] ),
    .S(_1639_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_1648_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5875_ (.A1(\as2650.stack_ptr[1] ),
    .A2(\as2650.stack_ptr[0] ),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5876_ (.I(_1649_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5877_ (.I(_1650_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5878_ (.A1(_1628_),
    .A2(_1651_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5879_ (.I(_1652_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5880_ (.I(_1653_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5881_ (.I(_1653_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5882_ (.A1(\as2650.stack[4][0] ),
    .A2(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5883_ (.A1(_1539_),
    .A2(_1654_),
    .B(_1656_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5884_ (.I(_1652_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5885_ (.I0(_1573_),
    .I1(\as2650.stack[4][1] ),
    .S(_1657_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5886_ (.I(_1658_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5887_ (.I0(_1579_),
    .I1(\as2650.stack[4][2] ),
    .S(_1657_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5888_ (.I(_1659_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_1653_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5890_ (.A1(\as2650.stack[4][3] ),
    .A2(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5891_ (.A1(_1583_),
    .A2(_1654_),
    .B(_1661_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5892_ (.I(_1653_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5893_ (.I0(_1589_),
    .I1(\as2650.stack[4][4] ),
    .S(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5894_ (.I(_1663_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(\as2650.stack[4][5] ),
    .A2(_1660_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5896_ (.A1(_1595_),
    .A2(_1654_),
    .B(_1664_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(\as2650.stack[4][6] ),
    .A2(_1660_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5898_ (.A1(_1600_),
    .A2(_1654_),
    .B(_1665_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5899_ (.A1(\as2650.stack[4][7] ),
    .A2(_1660_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5900_ (.A1(_1604_),
    .A2(_1655_),
    .B(_1666_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5901_ (.I0(_1610_),
    .I1(\as2650.stack[4][8] ),
    .S(_1662_),
    .Z(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1667_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5903_ (.A1(\as2650.stack[4][9] ),
    .A2(_1657_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5904_ (.A1(_1614_),
    .A2(_1655_),
    .B(_1668_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5905_ (.A1(\as2650.stack[4][10] ),
    .A2(_1657_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5906_ (.A1(_1617_),
    .A2(_1655_),
    .B(_1669_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5907_ (.I0(_1622_),
    .I1(\as2650.stack[4][11] ),
    .S(_1662_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_1670_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5909_ (.I0(_1626_),
    .I1(\as2650.stack[4][12] ),
    .S(_1662_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5910_ (.I(_1671_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5911_ (.I(_1536_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5912_ (.I(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5913_ (.I(\as2650.stack_ptr[1] ),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5914_ (.A1(_1541_),
    .A2(_1544_),
    .A3(_1564_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5915_ (.A1(_1674_),
    .A2(_1675_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5916_ (.I(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5917_ (.I0(\as2650.stack[1][0] ),
    .I1(_1673_),
    .S(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(_1678_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5919_ (.I(_1572_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5920_ (.I0(\as2650.stack[1][1] ),
    .I1(_1679_),
    .S(_1677_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5921_ (.I(_1680_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5922_ (.I(_1578_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5923_ (.I0(\as2650.stack[1][2] ),
    .I1(_1681_),
    .S(_1677_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5924_ (.I(_1682_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5925_ (.I(\as2650.pc[3] ),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5926_ (.I0(\as2650.stack[1][3] ),
    .I1(_1683_),
    .S(_1677_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_1684_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5928_ (.I(_1588_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5929_ (.I(_1676_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5930_ (.I0(\as2650.stack[1][4] ),
    .I1(_1685_),
    .S(_1686_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5931_ (.I(_1687_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5932_ (.I(\as2650.pc[5] ),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5933_ (.I(_1688_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5934_ (.I0(\as2650.stack[1][5] ),
    .I1(_1689_),
    .S(_1686_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5935_ (.I(_1690_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5936_ (.I(_1597_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5937_ (.I0(\as2650.stack[1][6] ),
    .I1(_1691_),
    .S(_1686_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5938_ (.I(_1692_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5939_ (.I(\as2650.pc[7] ),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5940_ (.I(_1693_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5941_ (.I0(\as2650.stack[1][7] ),
    .I1(_1694_),
    .S(_1686_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5942_ (.I(_1695_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5943_ (.I(_1609_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5944_ (.I(_1676_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5945_ (.I0(\as2650.stack[1][8] ),
    .I1(_1696_),
    .S(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5946_ (.I(_1698_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(\as2650.pc[9] ),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5948_ (.I(_1699_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5949_ (.I0(\as2650.stack[1][9] ),
    .I1(_1700_),
    .S(_1697_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_1701_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5951_ (.I(\as2650.pc[10] ),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5952_ (.I(_1702_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5953_ (.I0(\as2650.stack[1][10] ),
    .I1(_1703_),
    .S(_1697_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5954_ (.I(_1704_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5955_ (.I(_1621_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5956_ (.I0(\as2650.stack[1][11] ),
    .I1(_1705_),
    .S(_1697_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5957_ (.I(_1706_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5958_ (.I(_1625_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5959_ (.I0(\as2650.stack[1][12] ),
    .I1(_1707_),
    .S(_1676_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_1708_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5961_ (.I(_1538_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5962_ (.I(\as2650.stack_ptr[0] ),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5963_ (.I(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5964_ (.A1(\as2650.stack_ptr[1] ),
    .A2(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5965_ (.I(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5966_ (.I(_1713_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5967_ (.A1(_1628_),
    .A2(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5968_ (.I(_1715_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5969_ (.I(_1716_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_1716_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5971_ (.A1(\as2650.stack[5][0] ),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5972_ (.A1(_1709_),
    .A2(_1717_),
    .B(_1719_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5973_ (.I(_1715_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5974_ (.I0(_1573_),
    .I1(\as2650.stack[5][1] ),
    .S(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5975_ (.I(_1721_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5976_ (.I0(_1579_),
    .I1(\as2650.stack[5][2] ),
    .S(_1720_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5977_ (.I(_1722_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5978_ (.I(_1582_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5979_ (.I(_1716_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5980_ (.A1(\as2650.stack[5][3] ),
    .A2(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5981_ (.A1(_1723_),
    .A2(_1717_),
    .B(_1725_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5982_ (.I(_1716_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5983_ (.I0(_1589_),
    .I1(\as2650.stack[5][4] ),
    .S(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5984_ (.I(_1727_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5985_ (.A1(\as2650.stack[5][5] ),
    .A2(_1724_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5986_ (.A1(_1595_),
    .A2(_1717_),
    .B(_1728_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5987_ (.A1(\as2650.stack[5][6] ),
    .A2(_1724_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5988_ (.A1(_1600_),
    .A2(_1717_),
    .B(_1729_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5989_ (.A1(\as2650.stack[5][7] ),
    .A2(_1724_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5990_ (.A1(_1604_),
    .A2(_1718_),
    .B(_1730_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5991_ (.I0(_1610_),
    .I1(\as2650.stack[5][8] ),
    .S(_1726_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_1731_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5993_ (.I(_1613_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5994_ (.A1(\as2650.stack[5][9] ),
    .A2(_1720_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5995_ (.A1(_1732_),
    .A2(_1718_),
    .B(_1733_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_1616_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5997_ (.A1(\as2650.stack[5][10] ),
    .A2(_1720_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5998_ (.A1(_1734_),
    .A2(_1718_),
    .B(_1735_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5999_ (.I0(_1622_),
    .I1(\as2650.stack[5][11] ),
    .S(_1726_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_1736_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6001_ (.I0(_1626_),
    .I1(\as2650.stack[5][12] ),
    .S(_1726_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6002_ (.I(_1737_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6003_ (.A1(_1541_),
    .A2(_1564_),
    .A3(_1651_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6004_ (.I(_1738_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6005_ (.I(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6006_ (.I(_1739_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6007_ (.A1(\as2650.stack[0][0] ),
    .A2(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6008_ (.A1(_1709_),
    .A2(_1740_),
    .B(_1742_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6009_ (.I(_1738_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6010_ (.I0(_1679_),
    .I1(\as2650.stack[0][1] ),
    .S(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6011_ (.I(_1744_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6012_ (.I0(_1681_),
    .I1(\as2650.stack[0][2] ),
    .S(_1743_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6013_ (.I(_1745_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1739_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6015_ (.A1(\as2650.stack[0][3] ),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6016_ (.A1(_1723_),
    .A2(_1740_),
    .B(_1747_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6017_ (.I(_1739_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6018_ (.I0(_1685_),
    .I1(\as2650.stack[0][4] ),
    .S(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6019_ (.I(_1749_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6020_ (.A1(\as2650.stack[0][5] ),
    .A2(_1746_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6021_ (.A1(_1594_),
    .A2(_1740_),
    .B(_1750_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6022_ (.A1(\as2650.stack[0][6] ),
    .A2(_1746_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6023_ (.A1(_1599_),
    .A2(_1740_),
    .B(_1751_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6024_ (.A1(\as2650.stack[0][7] ),
    .A2(_1746_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6025_ (.A1(_1603_),
    .A2(_1741_),
    .B(_1752_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6026_ (.I0(_1696_),
    .I1(\as2650.stack[0][8] ),
    .S(_1748_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6027_ (.I(_1753_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6028_ (.A1(\as2650.stack[0][9] ),
    .A2(_1743_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6029_ (.A1(_1732_),
    .A2(_1741_),
    .B(_1754_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6030_ (.A1(\as2650.stack[0][10] ),
    .A2(_1743_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6031_ (.A1(_1734_),
    .A2(_1741_),
    .B(_1755_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6032_ (.I0(_1705_),
    .I1(\as2650.stack[0][11] ),
    .S(_1748_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6033_ (.I(_1756_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6034_ (.I0(_1707_),
    .I1(\as2650.stack[0][12] ),
    .S(_1748_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6035_ (.I(_1757_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6036_ (.A1(_1543_),
    .A2(_1675_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6037_ (.I(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6038_ (.I(_1759_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6039_ (.I(_1759_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(\as2650.stack[3][0] ),
    .A2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6041_ (.A1(_1709_),
    .A2(_1760_),
    .B(_1762_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6042_ (.I(_1758_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6043_ (.I0(_1679_),
    .I1(\as2650.stack[3][1] ),
    .S(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6044_ (.I(_1764_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6045_ (.I0(_1681_),
    .I1(\as2650.stack[3][2] ),
    .S(_1763_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6046_ (.I(_1765_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6047_ (.I(_1759_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6048_ (.A1(\as2650.stack[3][3] ),
    .A2(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6049_ (.A1(_1723_),
    .A2(_1760_),
    .B(_1767_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6050_ (.I(_1759_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6051_ (.I0(_1685_),
    .I1(\as2650.stack[3][4] ),
    .S(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6052_ (.I(_1769_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(\as2650.stack[3][5] ),
    .A2(_1766_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6054_ (.A1(_1594_),
    .A2(_1760_),
    .B(_1770_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6055_ (.A1(\as2650.stack[3][6] ),
    .A2(_1766_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6056_ (.A1(_1599_),
    .A2(_1760_),
    .B(_1771_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6057_ (.A1(\as2650.stack[3][7] ),
    .A2(_1766_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6058_ (.A1(_1603_),
    .A2(_1761_),
    .B(_1772_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6059_ (.I0(_1696_),
    .I1(\as2650.stack[3][8] ),
    .S(_1768_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_1773_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6061_ (.A1(\as2650.stack[3][9] ),
    .A2(_1763_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6062_ (.A1(_1732_),
    .A2(_1761_),
    .B(_1774_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6063_ (.A1(\as2650.stack[3][10] ),
    .A2(_1763_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6064_ (.A1(_1734_),
    .A2(_1761_),
    .B(_1775_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6065_ (.I0(_1705_),
    .I1(\as2650.stack[3][11] ),
    .S(_1768_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6066_ (.I(_1776_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6067_ (.I0(_1707_),
    .I1(\as2650.stack[3][12] ),
    .S(_1768_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_1777_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6069_ (.A1(_3848_),
    .A2(_1558_),
    .B(_1341_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6070_ (.A1(_0831_),
    .A2(_0938_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6071_ (.I(_1779_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6072_ (.A1(_1780_),
    .A2(_1252_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6073_ (.I(_1504_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6074_ (.I(_3548_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6075_ (.A1(_3771_),
    .A2(_1339_),
    .A3(_3524_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6076_ (.A1(_1244_),
    .A2(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6077_ (.I(_1785_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6078_ (.A1(_3545_),
    .A2(_1557_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6079_ (.I(_1787_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6080_ (.I(_1209_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6081_ (.A1(_1789_),
    .A2(_1340_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6082_ (.A1(_1783_),
    .A2(_1786_),
    .A3(_1788_),
    .A4(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6083_ (.A1(_1382_),
    .A2(_1782_),
    .A3(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6084_ (.I(\as2650.cycle[6] ),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6085_ (.I(_3601_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6086_ (.A1(_3586_),
    .A2(_1794_),
    .A3(_1238_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6087_ (.A1(_1793_),
    .A2(_1795_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6088_ (.A1(_3848_),
    .A2(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6089_ (.A1(_1778_),
    .A2(_1781_),
    .A3(_1792_),
    .A4(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6090_ (.A1(_3590_),
    .A2(_3602_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6091_ (.A1(_1793_),
    .A2(_1794_),
    .A3(_1238_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6092_ (.A1(_3586_),
    .A2(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6093_ (.A1(_1799_),
    .A2(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6094_ (.A1(_3586_),
    .A2(_1794_),
    .A3(_1239_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6095_ (.A1(_1558_),
    .A2(_1787_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6096_ (.A1(_1329_),
    .A2(_1803_),
    .A3(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6097_ (.A1(_1802_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6098_ (.A1(_1328_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6099_ (.I(_1788_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6100_ (.A1(_1331_),
    .A2(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_1783_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6102_ (.I(_1785_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6103_ (.I(_3674_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6104_ (.A1(_3514_),
    .A2(_1812_),
    .A3(_1782_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6105_ (.A1(_1810_),
    .A2(_1811_),
    .B(_1813_),
    .C(_1360_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6106_ (.I(_1265_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6107_ (.I(_1548_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6108_ (.I(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_1499_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_1498_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6111_ (.A1(_1815_),
    .A2(_1817_),
    .B(_1818_),
    .C(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6112_ (.A1(_3569_),
    .A2(_1784_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6113_ (.A1(_1498_),
    .A2(_1821_),
    .A3(_1554_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6114_ (.A1(_0311_),
    .A2(_1324_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6115_ (.A1(_1025_),
    .A2(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6116_ (.A1(_3547_),
    .A2(_1250_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6117_ (.A1(_1789_),
    .A2(_1785_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6118_ (.A1(_1783_),
    .A2(_1825_),
    .A3(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6119_ (.A1(_1820_),
    .A2(_1822_),
    .A3(_1824_),
    .A4(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6120_ (.A1(_1807_),
    .A2(_1809_),
    .A3(_1814_),
    .A4(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6121_ (.A1(_1798_),
    .A2(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6122_ (.I(_1830_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6123_ (.I(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6124_ (.I(\as2650.addr_buff[0] ),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6125_ (.I(_1830_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6126_ (.A1(_1833_),
    .A2(_1834_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6127_ (.A1(_1453_),
    .A2(_1832_),
    .B(_1835_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6128_ (.I(\as2650.addr_buff[1] ),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6129_ (.I(_1830_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6130_ (.A1(_1836_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6131_ (.A1(_1460_),
    .A2(_1832_),
    .B(_1838_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(\as2650.addr_buff[2] ),
    .A2(_1837_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6133_ (.A1(_0289_),
    .A2(_1832_),
    .B(_1839_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6134_ (.I(_1472_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6135_ (.I(\as2650.addr_buff[3] ),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6136_ (.A1(_1841_),
    .A2(_1837_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6137_ (.A1(_1840_),
    .A2(_1832_),
    .B(_1842_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6138_ (.I(_1480_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6139_ (.I(\as2650.addr_buff[4] ),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_1844_),
    .A2(_1837_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6141_ (.A1(_1843_),
    .A2(_1834_),
    .B(_1845_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6142_ (.I(_1483_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_3606_),
    .A2(_1831_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6144_ (.A1(_1846_),
    .A2(_1834_),
    .B(_1847_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6145_ (.I(_1456_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_3605_),
    .A2(_1831_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6147_ (.A1(_1848_),
    .A2(_1834_),
    .B(_1849_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6148_ (.I(_3846_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6149_ (.I0(_1525_),
    .I1(_1850_),
    .S(_1831_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_1851_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6151_ (.A1(_1210_),
    .A2(_1549_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6152_ (.I(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6153_ (.I(_1235_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_1854_),
    .A2(_1263_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6155_ (.A1(_1376_),
    .A2(_1246_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6156_ (.I(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6157_ (.A1(_1299_),
    .A2(_1855_),
    .A3(_1857_),
    .B(_1804_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6158_ (.A1(_3578_),
    .A2(_3570_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6159_ (.A1(_1854_),
    .A2(_1859_),
    .B(_1330_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6160_ (.I(_1248_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6161_ (.A1(_1853_),
    .A2(_1858_),
    .B(_1860_),
    .C(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6162_ (.A1(_1434_),
    .A2(_1322_),
    .B(_1809_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6163_ (.A1(net24),
    .A2(_1862_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6164_ (.A1(_1862_),
    .A2(_1863_),
    .B(_1864_),
    .C(_1280_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6165_ (.A1(_1241_),
    .A2(_1252_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6166_ (.A1(_3512_),
    .A2(_1235_),
    .A3(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6167_ (.A1(_1440_),
    .A2(_3570_),
    .A3(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6168_ (.A1(net22),
    .A2(_1867_),
    .B(_1431_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6169_ (.A1(_3770_),
    .A2(_1867_),
    .B(_1868_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6170_ (.I(net23),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6171_ (.I(_1342_),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6172_ (.I(_1870_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6173_ (.I(_1358_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6174_ (.I(_1872_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6175_ (.A1(_1375_),
    .A2(_1873_),
    .B(_1367_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_0939_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6177_ (.A1(_1875_),
    .A2(_1242_),
    .A3(_1859_),
    .A4(_1501_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6178_ (.I(_1789_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6179_ (.A1(_1877_),
    .A2(_1325_),
    .A3(_1859_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6180_ (.A1(_1254_),
    .A2(_1876_),
    .A3(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6181_ (.A1(_1871_),
    .A2(_1874_),
    .B(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6182_ (.A1(_3525_),
    .A2(_3526_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6183_ (.A1(_1881_),
    .A2(_1880_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6184_ (.I(_3513_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6185_ (.I(_1883_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6186_ (.A1(_1869_),
    .A2(_1880_),
    .B(_1882_),
    .C(_1884_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6187_ (.I(\as2650.cycle[7] ),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6188_ (.A1(_1885_),
    .A2(_3587_),
    .A3(_3588_),
    .A4(_3590_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6189_ (.A1(_3543_),
    .A2(_1240_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6190_ (.I(_1887_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6191_ (.A1(_1361_),
    .A2(_1232_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6192_ (.I(_1803_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6193_ (.A1(_1816_),
    .A2(_1889_),
    .A3(_1890_),
    .A4(_1804_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6194_ (.A1(_1888_),
    .A2(_1891_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6195_ (.A1(_1886_),
    .A2(_1806_),
    .A3(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6196_ (.A1(_1780_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6197_ (.A1(_1265_),
    .A2(_3536_),
    .A3(_1199_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6198_ (.I(_1784_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6199_ (.A1(_1819_),
    .A2(_1341_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6200_ (.I(_1897_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6201_ (.A1(_1253_),
    .A2(_1896_),
    .A3(_1898_),
    .B(_1272_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6202_ (.I(_3627_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6203_ (.A1(_1365_),
    .A2(_1900_),
    .B(_1335_),
    .C(_0359_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6204_ (.A1(_1309_),
    .A2(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6205_ (.A1(_1502_),
    .A2(_1897_),
    .B(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6206_ (.A1(_1895_),
    .A2(_1899_),
    .B(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(_1342_),
    .A2(_1362_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6208_ (.I(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6209_ (.A1(_1236_),
    .A2(_1905_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6210_ (.A1(_3581_),
    .A2(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6211_ (.A1(_1331_),
    .A2(_1808_),
    .B(_1878_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6212_ (.A1(_1505_),
    .A2(_1508_),
    .B(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6213_ (.A1(_1327_),
    .A2(_1906_),
    .B(_1908_),
    .C(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6214_ (.A1(_1366_),
    .A2(_1876_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6215_ (.A1(_1885_),
    .A2(_1800_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6216_ (.I(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6217_ (.A1(_1308_),
    .A2(_3600_),
    .A3(_1799_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6218_ (.A1(_1332_),
    .A2(_1914_),
    .B(_1915_),
    .C(_1360_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6219_ (.A1(_3496_),
    .A2(_3489_),
    .A3(_3535_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6220_ (.A1(_1216_),
    .A2(_1907_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_1793_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6222_ (.I(_1919_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6223_ (.I(_1890_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6224_ (.A1(_1920_),
    .A2(_1407_),
    .B(_1888_),
    .C(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6225_ (.A1(_1522_),
    .A2(_1917_),
    .A3(_1918_),
    .A4(_1922_),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6226_ (.A1(_1911_),
    .A2(_1912_),
    .A3(_1916_),
    .A4(_1923_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6227_ (.A1(_1894_),
    .A2(_1904_),
    .A3(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6228_ (.I(_1552_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6229_ (.A1(_3579_),
    .A2(_3692_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6230_ (.A1(_0284_),
    .A2(_0384_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6231_ (.A1(_3881_),
    .A2(_0494_),
    .A3(_1927_),
    .A4(_1928_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6232_ (.A1(_0576_),
    .A2(_0667_),
    .A3(_0780_),
    .A4(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_1197_),
    .A2(_1222_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6234_ (.A1(_0831_),
    .A2(_3779_),
    .A3(_1220_),
    .A4(_1221_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6235_ (.A1(_1931_),
    .A2(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6236_ (.A1(_1930_),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6237_ (.A1(_1528_),
    .A2(_1926_),
    .A3(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6238_ (.A1(_1925_),
    .A2(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6239_ (.I(_1871_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_1237_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6241_ (.I(_1938_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6242_ (.I(_3675_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6243_ (.I(_1940_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6244_ (.I(_3569_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6245_ (.A1(_1942_),
    .A2(_1818_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6246_ (.I(_1943_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6247_ (.I(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6248_ (.A1(_1250_),
    .A2(_1557_),
    .B(_0937_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6249_ (.A1(_1812_),
    .A2(_1941_),
    .B(_1945_),
    .C(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6250_ (.A1(net26),
    .A2(_1900_),
    .B(_1273_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6251_ (.A1(_1440_),
    .A2(_1939_),
    .A3(_1857_),
    .B1(_1947_),
    .B2(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6252_ (.A1(_1937_),
    .A2(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6253_ (.A1(net26),
    .A2(_1936_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6254_ (.A1(_1936_),
    .A2(_1950_),
    .B(_1951_),
    .C(_1280_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6255_ (.A1(_1526_),
    .A2(_1825_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6256_ (.I(_1352_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6257_ (.A1(_1953_),
    .A2(_1896_),
    .A3(_1550_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6258_ (.A1(_1386_),
    .A2(_1348_),
    .B(_1878_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6259_ (.A1(_1944_),
    .A2(_1952_),
    .B1(_1954_),
    .B2(_1332_),
    .C(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6260_ (.A1(_1318_),
    .A2(_1241_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6261_ (.A1(_1957_),
    .A2(_1501_),
    .A3(_1553_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_3671_),
    .A2(_3547_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6263_ (.A1(_3564_),
    .A2(_1959_),
    .B(_1943_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6264_ (.A1(_1958_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6265_ (.A1(_1263_),
    .A2(_1395_),
    .B(_1906_),
    .C(_1237_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6266_ (.A1(_1912_),
    .A2(_1961_),
    .A3(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6267_ (.A1(_1376_),
    .A2(_1908_),
    .B(_1956_),
    .C(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6268_ (.A1(_1903_),
    .A2(_1935_),
    .A3(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6269_ (.A1(net25),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6270_ (.I(_1446_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(_1783_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6272_ (.I(_1968_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6273_ (.I(_1969_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6274_ (.I(_1558_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6275_ (.A1(_1969_),
    .A2(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6276_ (.A1(_3846_),
    .A2(_1548_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6277_ (.I(_1973_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6278_ (.I(_1943_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6279_ (.A1(_1810_),
    .A2(_1975_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6280_ (.A1(_1553_),
    .A2(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6281_ (.A1(_1972_),
    .A2(_1974_),
    .B(_1977_),
    .C(_1780_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6282_ (.A1(_1812_),
    .A2(_1856_),
    .B1(_1946_),
    .B2(_1970_),
    .C(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6283_ (.A1(net25),
    .A2(_1526_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6284_ (.I(_0781_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6285_ (.A1(_1981_),
    .A2(_1504_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6286_ (.A1(_1979_),
    .A2(_1980_),
    .B(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6287_ (.A1(_1967_),
    .A2(_1983_),
    .B(_1522_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6288_ (.A1(_1937_),
    .A2(_1965_),
    .A3(_1984_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6289_ (.A1(_1280_),
    .A2(_1966_),
    .A3(_1985_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6290_ (.I(_1279_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6291_ (.I(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6292_ (.A1(_1373_),
    .A2(_1805_),
    .B(_1824_),
    .C(_1865_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6293_ (.A1(_1338_),
    .A2(_1891_),
    .A3(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6294_ (.I(_1241_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6295_ (.I(_1990_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6296_ (.A1(_1991_),
    .A2(_1989_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6297_ (.A1(_3555_),
    .A2(_1989_),
    .B1(_1992_),
    .B2(_3606_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6298_ (.A1(_1987_),
    .A2(_1993_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6299_ (.A1(_3554_),
    .A2(_1989_),
    .B1(_1992_),
    .B2(_3605_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6300_ (.A1(_1987_),
    .A2(_1994_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_1823_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6302_ (.I(_0698_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6303_ (.A1(_1365_),
    .A2(_0799_),
    .B1(_1995_),
    .B2(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(_1900_),
    .A2(_1901_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6305_ (.A1(_0698_),
    .A2(_1311_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6306_ (.I(_1266_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6307_ (.I(_2000_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6308_ (.A1(_0860_),
    .A2(_1362_),
    .A3(_1888_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6309_ (.A1(_1526_),
    .A2(_1335_),
    .B1(_1999_),
    .B2(_2001_),
    .C(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6310_ (.A1(_1997_),
    .A2(_1998_),
    .A3(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6311_ (.I(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6312_ (.I(_1267_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_0865_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6314_ (.A1(_1413_),
    .A2(_1439_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_2007_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6316_ (.A1(_2005_),
    .A2(_2009_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6317_ (.A1(_3759_),
    .A2(_2005_),
    .B(_2010_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6318_ (.I(_2006_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6319_ (.A1(_0908_),
    .A2(_2011_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6320_ (.A1(_1460_),
    .A2(_1307_),
    .B(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6321_ (.I0(_2013_),
    .I1(_3803_),
    .S(_2005_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6322_ (.I(_2014_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6323_ (.I(_1383_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6324_ (.I(_0280_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6325_ (.A1(_2016_),
    .A2(_1446_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6326_ (.A1(_0289_),
    .A2(_2015_),
    .B(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6327_ (.I0(_2018_),
    .I1(_3917_),
    .S(_2005_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6328_ (.I(_2019_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6329_ (.I(_0407_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6330_ (.A1(_2020_),
    .A2(_2011_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6331_ (.I(_1421_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6332_ (.I(_1272_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6333_ (.A1(_2022_),
    .A2(_2023_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2021_),
    .A2(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6335_ (.I(_2004_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6336_ (.I0(_2025_),
    .I1(_0339_),
    .S(_2026_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6337_ (.I(_2027_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6338_ (.I(_0492_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6339_ (.A1(_2028_),
    .A2(_2011_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6340_ (.A1(_1843_),
    .A2(_1307_),
    .B(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6341_ (.I0(_2030_),
    .I1(\as2650.holding_reg[4] ),
    .S(_2026_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6342_ (.I(_2031_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6343_ (.I(_1382_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6344_ (.A1(_1846_),
    .A2(_2032_),
    .B(_1268_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6345_ (.I0(_2033_),
    .I1(_0531_),
    .S(_2026_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6346_ (.I(_2034_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6347_ (.I(_2032_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6348_ (.I(_2035_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6349_ (.A1(_1425_),
    .A2(_1967_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6350_ (.A1(_1380_),
    .A2(_2036_),
    .B(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6351_ (.I0(_2038_),
    .I1(_0700_),
    .S(_2026_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6352_ (.I(_2039_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6353_ (.A1(_1525_),
    .A2(_1529_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6354_ (.A1(_1447_),
    .A2(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6355_ (.I0(_2041_),
    .I1(_0737_),
    .S(_2004_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6356_ (.I(_2042_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6357_ (.A1(_2036_),
    .A2(_1334_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6358_ (.I(_3519_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6359_ (.I(_2044_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6360_ (.A1(_1338_),
    .A2(_2043_),
    .B(_2045_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6361_ (.I(_1248_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6362_ (.I(\as2650.cycle[0] ),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6363_ (.I(_1782_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6365_ (.A1(_2047_),
    .A2(_1382_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6366_ (.I(_1217_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6367_ (.I(_3581_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6368_ (.I(_3611_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6369_ (.A1(_2051_),
    .A2(_1223_),
    .B(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6370_ (.A1(_2051_),
    .A2(_2052_),
    .A3(_1895_),
    .B(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6371_ (.I(_1816_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6372_ (.I(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6373_ (.A1(_2057_),
    .A2(_1326_),
    .A3(_1859_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6374_ (.I(_1817_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6375_ (.I(_1786_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6376_ (.A1(_1850_),
    .A2(_2059_),
    .B1(_1959_),
    .B2(_3526_),
    .C(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6377_ (.A1(_1385_),
    .A2(_1930_),
    .A3(_1933_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6378_ (.A1(_1969_),
    .A2(_2050_),
    .B(_2062_),
    .C(_1944_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6379_ (.A1(_2061_),
    .A2(_2063_),
    .B(_1553_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6380_ (.A1(_2050_),
    .A2(_2055_),
    .B(_2058_),
    .C(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6381_ (.A1(_2047_),
    .A2(_2049_),
    .B1(_1865_),
    .B2(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6382_ (.A1(_1320_),
    .A2(_2066_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6383_ (.I(_1373_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6384_ (.I(_0315_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6385_ (.I(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6386_ (.I(_3876_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_1886_),
    .A2(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6388_ (.A1(_3526_),
    .A2(_1886_),
    .B(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6389_ (.I(_0940_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6390_ (.I(_1799_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6391_ (.A1(_1850_),
    .A2(_2071_),
    .B(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6392_ (.A1(_1919_),
    .A2(_1795_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6393_ (.I(_2077_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6394_ (.A1(_1407_),
    .A2(_2071_),
    .B(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6395_ (.A1(_1439_),
    .A2(_2074_),
    .A3(_2076_),
    .A4(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6396_ (.A1(_2070_),
    .A2(_2073_),
    .B(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_1323_),
    .A2(_1465_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6398_ (.A1(_2068_),
    .A2(_1906_),
    .A3(_2081_),
    .A4(_2082_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6399_ (.A1(_2067_),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6400_ (.A1(_2046_),
    .A2(_2047_),
    .B1(_1254_),
    .B2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6401_ (.A1(_1987_),
    .A2(_2085_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6402_ (.I(_1861_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6403_ (.A1(_2086_),
    .A2(_3525_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6404_ (.A1(_2000_),
    .A2(_1934_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6405_ (.A1(_3525_),
    .A2(_2047_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6406_ (.I(_1818_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(_1272_),
    .A2(_1971_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6408_ (.A1(_2090_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6409_ (.A1(_2089_),
    .A2(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6410_ (.A1(_1881_),
    .A2(_1959_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6411_ (.A1(_1521_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6412_ (.A1(_2089_),
    .A2(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6413_ (.A1(_2088_),
    .A2(_2093_),
    .B1(_2096_),
    .B2(_1896_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6414_ (.A1(_1338_),
    .A2(_1342_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6415_ (.I(_1796_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6416_ (.A1(_2072_),
    .A2(_2076_),
    .A3(_2089_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6417_ (.A1(_2099_),
    .A2(_2100_),
    .B(_2091_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6418_ (.A1(_2079_),
    .A2(_2101_),
    .B(_2082_),
    .C(_1433_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6419_ (.A1(_1273_),
    .A2(_2089_),
    .B(_2055_),
    .C(_1320_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6420_ (.A1(_2098_),
    .A2(_2102_),
    .A3(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6421_ (.A1(_1340_),
    .A2(_2097_),
    .B(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6422_ (.A1(_2087_),
    .A2(_2105_),
    .B(_2045_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6423_ (.I(_2053_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6424_ (.I(_2106_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6425_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6426_ (.I(_3564_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6427_ (.A1(_1556_),
    .A2(_2109_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6428_ (.A1(_1527_),
    .A2(_2052_),
    .B1(_1853_),
    .B2(_1857_),
    .C(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6429_ (.I(_1217_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6430_ (.I(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6431_ (.A1(_3672_),
    .A2(_2109_),
    .A3(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6432_ (.A1(_1527_),
    .A2(_1857_),
    .B(_2111_),
    .C(_2114_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6433_ (.I(_2106_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6434_ (.A1(_1527_),
    .A2(_2049_),
    .A3(_2110_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6435_ (.I(_1968_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6436_ (.A1(_2118_),
    .A2(_2110_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6437_ (.A1(_2094_),
    .A2(_2119_),
    .B(_1974_),
    .C(_1945_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6438_ (.I(_1811_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6439_ (.A1(_2121_),
    .A2(_2119_),
    .B(_2048_),
    .C(_1554_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6440_ (.A1(_2120_),
    .A2(_2122_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6441_ (.A1(_2116_),
    .A2(_2117_),
    .A3(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6442_ (.I(_1957_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_2125_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6444_ (.I(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6445_ (.A1(_2108_),
    .A2(_2115_),
    .B(_2124_),
    .C(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6446_ (.A1(_1996_),
    .A2(_1336_),
    .B(_2119_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6447_ (.A1(_1888_),
    .A2(_2129_),
    .B(_2046_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6448_ (.I(_1279_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6449_ (.A1(_2086_),
    .A2(_3546_),
    .B1(_2128_),
    .B2(_2130_),
    .C(_2131_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6450_ (.I(_1279_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6451_ (.A1(\as2650.cycle[3] ),
    .A2(_1556_),
    .A3(_2109_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6452_ (.A1(_1556_),
    .A2(_2109_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6453_ (.A1(_1555_),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6454_ (.A1(_2133_),
    .A2(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_2078_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6456_ (.A1(_1448_),
    .A2(_2077_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6457_ (.A1(_0973_),
    .A2(_2137_),
    .B(_2138_),
    .C(_2071_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6458_ (.A1(_2072_),
    .A2(_2136_),
    .A3(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6459_ (.A1(_1970_),
    .A2(_1971_),
    .B(_1926_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6460_ (.A1(_1408_),
    .A2(_1322_),
    .A3(_2049_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6461_ (.A1(_1926_),
    .A2(_1974_),
    .B1(_2136_),
    .B2(_2141_),
    .C(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6462_ (.A1(_1946_),
    .A2(_2140_),
    .B1(_2143_),
    .B2(_1442_),
    .C(_1861_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6463_ (.A1(_2086_),
    .A2(_1555_),
    .B(_2132_),
    .C(_2144_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6464_ (.I(_3588_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6465_ (.A1(_1248_),
    .A2(_2133_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6466_ (.A1(_2145_),
    .A2(_2146_),
    .B(_1431_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6467_ (.A1(_2145_),
    .A2(_2146_),
    .B(_2147_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6468_ (.A1(_2145_),
    .A2(_2146_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6469_ (.A1(_3587_),
    .A2(_2148_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6470_ (.A1(_1987_),
    .A2(_2149_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6471_ (.A1(_1920_),
    .A2(_1884_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6472_ (.A1(_1320_),
    .A2(_1871_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(_3587_),
    .A2(_2145_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6474_ (.A1(_2133_),
    .A2(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6475_ (.A1(_1920_),
    .A2(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6476_ (.A1(_3591_),
    .A2(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6477_ (.A1(_0973_),
    .A2(_2155_),
    .B(_2138_),
    .C(_1440_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6478_ (.A1(_1307_),
    .A2(_1550_),
    .B(_2151_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6479_ (.A1(_2151_),
    .A2(_2154_),
    .B1(_2156_),
    .B2(_2157_),
    .C(_2046_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6480_ (.A1(_1503_),
    .A2(_2150_),
    .B(_2158_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6481_ (.I(_1430_),
    .Z(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6482_ (.A1(_1885_),
    .A2(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6483_ (.I(_1995_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6484_ (.I(_2161_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6485_ (.A1(_1920_),
    .A2(_2153_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6486_ (.A1(_1885_),
    .A2(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6487_ (.A1(_1025_),
    .A2(_2162_),
    .A3(_1797_),
    .A4(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6488_ (.A1(_2108_),
    .A2(_2162_),
    .B(_2165_),
    .C(_2046_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6489_ (.A1(_1503_),
    .A2(_2160_),
    .B(_2166_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6490_ (.A1(_1793_),
    .A2(_1890_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6491_ (.A1(_0831_),
    .A2(_1913_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6492_ (.A1(_3611_),
    .A2(_3576_),
    .B(_1915_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6493_ (.A1(_1778_),
    .A2(_2168_),
    .A3(_2169_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6494_ (.A1(_3591_),
    .A2(_1807_),
    .B1(_2167_),
    .B2(_1330_),
    .C(_2170_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6495_ (.A1(_1900_),
    .A2(_1808_),
    .A3(_2138_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6496_ (.A1(_3570_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_3676_),
    .A2(_1360_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6498_ (.A1(_1318_),
    .A2(_1326_),
    .B1(_1856_),
    .B2(_1815_),
    .C(_0860_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6499_ (.A1(_1995_),
    .A2(_1781_),
    .A3(_2174_),
    .A4(_2175_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6500_ (.A1(_2171_),
    .A2(_2173_),
    .A3(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6501_ (.I(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6502_ (.I(_2178_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6503_ (.I(_0974_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6504_ (.I(_2180_),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6505_ (.I(_0974_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6506_ (.A1(_2182_),
    .A2(_0883_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6507_ (.A1(_0865_),
    .A2(_2181_),
    .B(_2183_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6508_ (.I(_2177_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(net41),
    .A2(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6510_ (.A1(_2179_),
    .A2(_2184_),
    .B(_2186_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6511_ (.I(_0974_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6512_ (.I(_3816_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6513_ (.I(_0908_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6514_ (.A1(_2189_),
    .A2(_2187_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6515_ (.A1(_2187_),
    .A2(_2188_),
    .B(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6516_ (.I(_2177_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6517_ (.A1(net42),
    .A2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6518_ (.A1(_2179_),
    .A2(_2191_),
    .B(_2193_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6519_ (.A1(_2182_),
    .A2(_0960_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6520_ (.A1(_2016_),
    .A2(_2181_),
    .B(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6521_ (.A1(net43),
    .A2(_2192_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6522_ (.A1(_2179_),
    .A2(_2195_),
    .B(_2196_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6523_ (.I(_0307_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6524_ (.I0(_2197_),
    .I1(_2020_),
    .S(_2180_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6525_ (.I0(_2198_),
    .I1(net44),
    .S(_2178_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6526_ (.I(_2199_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6527_ (.A1(_2180_),
    .A2(_0561_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6528_ (.A1(_2028_),
    .A2(_2181_),
    .B(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6529_ (.A1(net45),
    .A2(_2192_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6530_ (.A1(_2179_),
    .A2(_2201_),
    .B(_2202_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6531_ (.A1(_2180_),
    .A2(_1096_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6532_ (.A1(_1017_),
    .A2(_2181_),
    .B(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6533_ (.A1(net19),
    .A2(_2192_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6534_ (.A1(_2185_),
    .A2(_2204_),
    .B(_2205_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6535_ (.A1(_1380_),
    .A2(_2182_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6536_ (.A1(_2187_),
    .A2(_0706_),
    .B(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(net20),
    .A2(_2178_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6538_ (.A1(_2185_),
    .A2(_2207_),
    .B(_2208_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6539_ (.A1(_1114_),
    .A2(_2182_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6540_ (.A1(_2187_),
    .A2(_1101_),
    .B(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6541_ (.A1(net21),
    .A2(_2178_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6542_ (.A1(_2185_),
    .A2(_2210_),
    .B(_2211_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6543_ (.I(net4),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6544_ (.A1(_2212_),
    .A2(_1196_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6545_ (.I(_2015_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6546_ (.A1(_1113_),
    .A2(_1196_),
    .B(_2213_),
    .C(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6547_ (.I(_1448_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_1159_),
    .A2(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6549_ (.A1(\as2650.psu[7] ),
    .A2(_1408_),
    .B(_1353_),
    .C(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6550_ (.A1(_2212_),
    .A2(_1353_),
    .B(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6551_ (.A1(_1529_),
    .A2(_2219_),
    .B(_1861_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6552_ (.A1(_1481_),
    .A2(_2086_),
    .B1(_2215_),
    .B2(_2220_),
    .C(_2131_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6553_ (.A1(_3543_),
    .A2(_1355_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6554_ (.A1(_1246_),
    .A2(_1216_),
    .A3(_1356_),
    .A4(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6555_ (.A1(_1887_),
    .A2(_1804_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6556_ (.A1(_1359_),
    .A2(_1366_),
    .A3(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6557_ (.A1(_2222_),
    .A2(_1865_),
    .B(_1903_),
    .C(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6558_ (.A1(_0939_),
    .A2(_1971_),
    .A3(_1786_),
    .A4(_1788_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6559_ (.A1(_1958_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6560_ (.A1(_1197_),
    .A2(_1222_),
    .A3(_2082_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6561_ (.A1(_0312_),
    .A2(_1796_),
    .B(_2228_),
    .C(_3511_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6562_ (.A1(_1788_),
    .A2(_1973_),
    .B(_1552_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6563_ (.A1(_0311_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6564_ (.A1(_1811_),
    .A2(_1974_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6565_ (.A1(_1961_),
    .A2(_2227_),
    .A3(_2229_),
    .A4(_2232_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6566_ (.A1(_1324_),
    .A2(_1216_),
    .A3(_1907_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6567_ (.A1(_1361_),
    .A2(_1917_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6568_ (.A1(_1367_),
    .A2(_1341_),
    .B(_2235_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6569_ (.A1(_1210_),
    .A2(_1786_),
    .A3(_1825_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6570_ (.A1(_1351_),
    .A2(_1982_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6571_ (.A1(_1779_),
    .A2(_1226_),
    .A3(_2237_),
    .A4(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6572_ (.A1(_1908_),
    .A2(_2234_),
    .A3(_2236_),
    .A4(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6573_ (.A1(_1892_),
    .A2(_2225_),
    .A3(_2233_),
    .A4(_2240_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6574_ (.I(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6575_ (.I(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6576_ (.I(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6577_ (.I(_1821_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6578_ (.I(_2245_),
    .Z(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6579_ (.A1(_1872_),
    .A2(_1944_),
    .B(_2062_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6580_ (.I(_1519_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6581_ (.A1(_1538_),
    .A2(_2248_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6582_ (.A1(_1385_),
    .A2(_1934_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6583_ (.A1(_2060_),
    .A2(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6584_ (.I(\as2650.addr_buff[0] ),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6585_ (.I(_2252_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6586_ (.A1(_1536_),
    .A2(_3665_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6587_ (.A1(_1537_),
    .A2(_1519_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6588_ (.A1(_1519_),
    .A2(_2254_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6589_ (.A1(_3666_),
    .A2(_0939_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6590_ (.A1(_2253_),
    .A2(_1852_),
    .B1(_2256_),
    .B2(_1877_),
    .C(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6591_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_3481_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(_1816_),
    .A2(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6593_ (.A1(_3667_),
    .A2(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6594_ (.A1(_1412_),
    .A2(_2260_),
    .B(_2261_),
    .C(_1826_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6595_ (.A1(_1975_),
    .A2(_2258_),
    .B(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6596_ (.A1(_1386_),
    .A2(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6597_ (.A1(_1538_),
    .A2(_2247_),
    .B1(_2249_),
    .B2(_2251_),
    .C(_2264_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6598_ (.A1(_1438_),
    .A2(_2245_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_1438_),
    .A2(_1782_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6600_ (.A1(_2254_),
    .A2(_2267_),
    .B(_2106_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6601_ (.A1(_2246_),
    .A2(_2265_),
    .B1(_2266_),
    .B2(_1672_),
    .C(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6602_ (.A1(\as2650.stack_ptr[2] ),
    .A2(_1649_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6603_ (.I(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6604_ (.I(_1712_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6605_ (.A1(_1542_),
    .A2(_1710_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(_2273_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6607_ (.I(_2274_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6608_ (.A1(\as2650.stack[4][0] ),
    .A2(_2272_),
    .B1(_2275_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6609_ (.I(_1546_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_1650_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6611_ (.A1(\as2650.stack[5][0] ),
    .A2(_2277_),
    .B1(_2278_),
    .B2(\as2650.stack[7][0] ),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6612_ (.A1(_2271_),
    .A2(_2276_),
    .A3(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6613_ (.A1(_1540_),
    .A2(_1649_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6614_ (.I(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(_1649_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_2273_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6617_ (.A1(\as2650.stack[3][0] ),
    .A2(_2283_),
    .B1(_2284_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6618_ (.I(_1545_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6619_ (.I(_1712_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6620_ (.A1(\as2650.stack[1][0] ),
    .A2(_2286_),
    .B1(_2287_),
    .B2(\as2650.stack[0][0] ),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6621_ (.A1(_2282_),
    .A2(_2285_),
    .A3(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6622_ (.A1(_2280_),
    .A2(_2289_),
    .B(_1204_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6623_ (.A1(_1672_),
    .A2(_1264_),
    .B(_2290_),
    .C(_2116_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6624_ (.A1(_2269_),
    .A2(_2291_),
    .B(_2126_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6625_ (.I(_2241_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6626_ (.A1(_1673_),
    .A2(_2127_),
    .B(_2292_),
    .C(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6627_ (.A1(_1884_),
    .A2(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6628_ (.A1(_1539_),
    .A2(_2244_),
    .B(_2295_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6629_ (.I(_1986_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6630_ (.I(_2241_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6631_ (.I(_2297_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6632_ (.A1(_1570_),
    .A2(_1536_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6633_ (.I(_2299_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6634_ (.A1(\as2650.pc[0] ),
    .A2(net5),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6635_ (.A1(\as2650.pc[1] ),
    .A2(net6),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6636_ (.A1(_2301_),
    .A2(_2302_),
    .Z(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6637_ (.I(_1821_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6638_ (.A1(_1815_),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6639_ (.I(_2305_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6640_ (.A1(_1930_),
    .A2(_1933_),
    .B(_1815_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6641_ (.I(_2307_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6642_ (.I(_1206_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6643_ (.A1(_1537_),
    .A2(_2309_),
    .B(_1571_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6644_ (.A1(_1571_),
    .A2(_1672_),
    .A3(_2309_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6645_ (.A1(_2310_),
    .A2(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6646_ (.I(\as2650.addr_buff[1] ),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6647_ (.I(_2313_),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6648_ (.A1(_0894_),
    .A2(_1549_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6649_ (.A1(_2314_),
    .A2(_2056_),
    .B(_2315_),
    .C(_1352_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6650_ (.A1(_1942_),
    .A2(_2303_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6651_ (.A1(_2309_),
    .A2(_2299_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6652_ (.A1(_1211_),
    .A2(_2317_),
    .A3(_2318_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6653_ (.A1(_1438_),
    .A2(_2316_),
    .A3(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6654_ (.A1(_2308_),
    .A2(_2312_),
    .B(_2320_),
    .C(_2060_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6655_ (.A1(_2062_),
    .A2(_2299_),
    .B(_2321_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6656_ (.A1(_1872_),
    .A2(_1975_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6657_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_0396_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6658_ (.A1(_3882_),
    .A2(_2324_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6659_ (.A1(_1412_),
    .A2(_2259_),
    .B(_2325_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_1817_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6661_ (.A1(net5),
    .A2(_2259_),
    .A3(_2325_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_2327_),
    .A2(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6663_ (.A1(_1415_),
    .A2(_1875_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6664_ (.A1(_1358_),
    .A2(_1811_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6665_ (.A1(_2326_),
    .A2(_2329_),
    .B(_2330_),
    .C(_2331_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6666_ (.I(_2245_),
    .Z(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6667_ (.A1(_2323_),
    .A2(_2300_),
    .B(_2332_),
    .C(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6668_ (.A1(_2322_),
    .A2(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6669_ (.A1(_2266_),
    .A2(_2300_),
    .B1(_2303_),
    .B2(_2306_),
    .C(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6670_ (.A1(_0937_),
    .A2(_1870_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6671_ (.I(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6672_ (.I(_2051_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6673_ (.I(_1546_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6674_ (.A1(\as2650.stack[5][1] ),
    .A2(_2340_),
    .B1(_1714_),
    .B2(\as2650.stack[4][1] ),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6675_ (.I(_1650_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_2274_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6677_ (.A1(\as2650.stack[7][1] ),
    .A2(_2342_),
    .B1(_2343_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6678_ (.A1(_2271_),
    .A2(_2341_),
    .A3(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_2281_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6680_ (.A1(\as2650.stack[1][1] ),
    .A2(_1547_),
    .B1(_1714_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6681_ (.A1(\as2650.stack[3][1] ),
    .A2(_2342_),
    .B1(_2343_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6682_ (.A1(_2346_),
    .A2(_2347_),
    .A3(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6683_ (.A1(_2339_),
    .A2(_2345_),
    .A3(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6684_ (.A1(_1204_),
    .A2(_2300_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6685_ (.A1(_2350_),
    .A2(_2351_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_1243_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6687_ (.A1(_2338_),
    .A2(_2300_),
    .B1(_2352_),
    .B2(_2353_),
    .C(_2242_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6688_ (.A1(_1898_),
    .A2(_2336_),
    .B(_2354_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6689_ (.A1(_1572_),
    .A2(_2298_),
    .B(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6690_ (.A1(_2296_),
    .A2(_2356_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6691_ (.I(_2297_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6692_ (.A1(_1578_),
    .A2(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_2242_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6694_ (.A1(_1570_),
    .A2(_1537_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6695_ (.A1(_1577_),
    .A2(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6696_ (.I(_2247_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6697_ (.A1(_2000_),
    .A2(_1505_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6698_ (.I(_2363_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6699_ (.I(_1942_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6700_ (.A1(\as2650.pc[1] ),
    .A2(_3882_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6701_ (.A1(_2301_),
    .A2(_2302_),
    .B(_2366_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6702_ (.A1(\as2650.pc[2] ),
    .A2(net7),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6703_ (.A1(_2367_),
    .A2(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6704_ (.A1(_2367_),
    .A2(_2368_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6705_ (.A1(_2365_),
    .A2(_2369_),
    .A3(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6706_ (.A1(_1383_),
    .A2(_2090_),
    .A3(_2371_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6707_ (.I(_2106_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6708_ (.A1(_2364_),
    .A2(_2361_),
    .B(_2372_),
    .C(_2373_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6709_ (.I(_2125_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6710_ (.A1(_2362_),
    .A2(_2374_),
    .B(_2375_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6711_ (.I(_2060_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6712_ (.I(_2307_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6713_ (.A1(_1577_),
    .A2(_2310_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6714_ (.I(_1942_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6715_ (.I(_1877_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6716_ (.A1(_2380_),
    .A2(_2361_),
    .B(_2371_),
    .C(_2381_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6717_ (.I(\as2650.addr_buff[2] ),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6718_ (.I(_2056_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6719_ (.I(_1549_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6720_ (.A1(_1417_),
    .A2(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6721_ (.A1(_2383_),
    .A2(_2384_),
    .B(_1233_),
    .C(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6722_ (.A1(_2378_),
    .A2(_2379_),
    .B(_2382_),
    .C(_2387_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6723_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_3480_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6724_ (.A1(_0285_),
    .A2(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6725_ (.A1(_0285_),
    .A2(_2389_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6726_ (.A1(_3883_),
    .A2(_2324_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6727_ (.A1(_2390_),
    .A2(_2391_),
    .B(_2392_),
    .C(_2328_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _6728_ (.A1(_2392_),
    .A2(_2328_),
    .B(_2390_),
    .C(_2391_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6729_ (.A1(_2118_),
    .A2(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6730_ (.A1(_1418_),
    .A2(_1875_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6731_ (.A1(_2331_),
    .A2(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6732_ (.A1(_2393_),
    .A2(_2395_),
    .B(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6733_ (.A1(_2377_),
    .A2(_2388_),
    .B(_2398_),
    .C(_2049_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_2274_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6735_ (.A1(\as2650.stack[7][2] ),
    .A2(_2342_),
    .B1(_2400_),
    .B2(\as2650.stack[6][2] ),
    .C1(_1714_),
    .C2(\as2650.stack[4][2] ),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6736_ (.I(_2286_),
    .Z(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6737_ (.A1(\as2650.stack[5][2] ),
    .A2(_2402_),
    .B(_2346_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6738_ (.A1(\as2650.stack[1][2] ),
    .A2(_2286_),
    .B1(_1713_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6739_ (.A1(_2282_),
    .A2(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6740_ (.A1(\as2650.stack[3][2] ),
    .A2(_1651_),
    .B1(_2400_),
    .B2(\as2650.stack[2][2] ),
    .C(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6741_ (.A1(_2401_),
    .A2(_2403_),
    .B(_2406_),
    .C(_1264_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6742_ (.I(_2051_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6743_ (.I(_1854_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6744_ (.A1(_2408_),
    .A2(_2361_),
    .B(_2409_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6745_ (.A1(_2374_),
    .A2(_2399_),
    .B1(_2407_),
    .B2(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6746_ (.A1(_2361_),
    .A2(_2376_),
    .B1(_2411_),
    .B2(_2127_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6747_ (.A1(_2359_),
    .A2(_2412_),
    .B(_2159_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6748_ (.A1(_2358_),
    .A2(_2413_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6749_ (.A1(_1576_),
    .A2(\as2650.pc[1] ),
    .A3(_1535_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6750_ (.A1(_1683_),
    .A2(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6751_ (.A1(\as2650.pc[3] ),
    .A2(net8),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6752_ (.A1(_1581_),
    .A2(_1471_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6753_ (.A1(_2416_),
    .A2(_2417_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6754_ (.A1(_1576_),
    .A2(_0285_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6755_ (.A1(_2419_),
    .A2(_2370_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6756_ (.A1(_2418_),
    .A2(_2420_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6757_ (.I(_2267_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6758_ (.A1(_2364_),
    .A2(_2415_),
    .B1(_2421_),
    .B2(_2422_),
    .C(_2373_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6759_ (.A1(_2362_),
    .A2(_2423_),
    .B(_2375_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6760_ (.A1(_1535_),
    .A2(_3573_),
    .B(_1576_),
    .C(_1570_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6761_ (.A1(_1582_),
    .A2(_2425_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6762_ (.I(_1968_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6763_ (.A1(_1841_),
    .A2(_1875_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6764_ (.A1(_1840_),
    .A2(_2427_),
    .B(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6765_ (.I(_2309_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6766_ (.A1(_2365_),
    .A2(_2415_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6767_ (.A1(_2430_),
    .A2(_2421_),
    .B(_2431_),
    .C(_2381_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6768_ (.A1(_2308_),
    .A2(_2426_),
    .B1(_2429_),
    .B2(_1873_),
    .C(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6769_ (.I(_2331_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6770_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_3481_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6771_ (.A1(net8),
    .A2(_2435_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6772_ (.A1(_2390_),
    .A2(_2394_),
    .A3(_2436_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6773_ (.A1(_2390_),
    .A2(_2394_),
    .B(_2436_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6774_ (.A1(_2384_),
    .A2(_2437_),
    .A3(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6775_ (.A1(_1420_),
    .A2(_1969_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6776_ (.A1(_2434_),
    .A2(_2439_),
    .A3(_2440_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6777_ (.I(_1505_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6778_ (.A1(_2377_),
    .A2(_2433_),
    .B(_2441_),
    .C(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6779_ (.I(_2270_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6780_ (.I(_1650_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6781_ (.A1(\as2650.stack[5][3] ),
    .A2(_2277_),
    .B1(_2445_),
    .B2(\as2650.stack[7][3] ),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6782_ (.I(_1712_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6783_ (.I(_2274_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6784_ (.A1(\as2650.stack[4][3] ),
    .A2(_2447_),
    .B1(_2448_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6785_ (.A1(_2444_),
    .A2(_2446_),
    .A3(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6786_ (.I(_1546_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6787_ (.A1(\as2650.stack[1][3] ),
    .A2(_2451_),
    .B1(_2275_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6788_ (.A1(\as2650.stack[3][3] ),
    .A2(_2445_),
    .B1(_2287_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6789_ (.A1(_2282_),
    .A2(_2452_),
    .A3(_2453_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6790_ (.A1(_1218_),
    .A2(_2450_),
    .A3(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6791_ (.I(_1854_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6792_ (.A1(_2408_),
    .A2(_2415_),
    .B(_2455_),
    .C(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6793_ (.A1(_2423_),
    .A2(_2443_),
    .B(_2457_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6794_ (.I(_2126_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6795_ (.A1(_2415_),
    .A2(_2424_),
    .B1(_2458_),
    .B2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6796_ (.I(_1430_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6797_ (.A1(_2243_),
    .A2(_2460_),
    .B(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6798_ (.A1(_1583_),
    .A2(_2244_),
    .B(_2462_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6799_ (.A1(_1588_),
    .A2(_2359_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6800_ (.I(_2363_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6801_ (.A1(_1581_),
    .A2(_2414_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6802_ (.A1(_1586_),
    .A2(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6804_ (.A1(\as2650.pc[4] ),
    .A2(_1477_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6805_ (.I(_2416_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6806_ (.A1(_2469_),
    .A2(_2420_),
    .B(_2417_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6807_ (.A1(_2468_),
    .A2(_2470_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6808_ (.A1(_2306_),
    .A2(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6809_ (.I(_2053_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6810_ (.I(_2473_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6811_ (.I(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6812_ (.A1(_2464_),
    .A2(_2467_),
    .B(_2472_),
    .C(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6813_ (.A1(_2088_),
    .A2(_2323_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6814_ (.I(_2477_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6815_ (.I(_2333_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6816_ (.A1(_1581_),
    .A2(_2425_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6817_ (.A1(_1587_),
    .A2(_2480_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6818_ (.I(\as2650.addr_buff[4] ),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6819_ (.A1(_2365_),
    .A2(_2466_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6820_ (.A1(_2380_),
    .A2(_2471_),
    .B(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6821_ (.A1(_1423_),
    .A2(_1810_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6822_ (.A1(_2482_),
    .A2(_1852_),
    .B1(_2484_),
    .B2(_2381_),
    .C(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6823_ (.A1(_2378_),
    .A2(_2481_),
    .B1(_2486_),
    .B2(_2006_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6824_ (.A1(_0386_),
    .A2(_2435_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6825_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_3481_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6826_ (.A1(net9),
    .A2(_2489_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6827_ (.I(_2490_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6828_ (.A1(_2488_),
    .A2(_2438_),
    .A3(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6829_ (.I(_1810_),
    .Z(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6830_ (.A1(_2488_),
    .A2(_2438_),
    .B(_2491_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6831_ (.A1(_2493_),
    .A2(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6832_ (.A1(_2492_),
    .A2(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6833_ (.A1(_1232_),
    .A2(_1975_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6834_ (.I(_2497_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6835_ (.A1(_1479_),
    .A2(_1817_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6836_ (.A1(_2498_),
    .A2(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6837_ (.A1(_2090_),
    .A2(_2487_),
    .B1(_2496_),
    .B2(_2500_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6838_ (.A1(_2479_),
    .A2(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6839_ (.I(_2125_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6840_ (.A1(_2478_),
    .A2(_2467_),
    .B1(_2502_),
    .B2(_2503_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6841_ (.I(_2112_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6842_ (.I(_2282_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6843_ (.I(_2283_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6844_ (.I(_2287_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6845_ (.A1(\as2650.stack[3][4] ),
    .A2(_2507_),
    .B1(_2508_),
    .B2(\as2650.stack[0][4] ),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6846_ (.I(_2284_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6847_ (.A1(\as2650.stack[1][4] ),
    .A2(_2402_),
    .B1(_2510_),
    .B2(\as2650.stack[2][4] ),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6848_ (.A1(_2506_),
    .A2(_2509_),
    .A3(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6849_ (.I(_2270_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6850_ (.A1(\as2650.stack[5][4] ),
    .A2(_2402_),
    .B1(_2510_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6851_ (.A1(\as2650.stack[7][4] ),
    .A2(_2507_),
    .B1(_2508_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6852_ (.A1(_2513_),
    .A2(_2514_),
    .A3(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6853_ (.A1(_2505_),
    .A2(_2512_),
    .A3(_2516_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6854_ (.A1(_2113_),
    .A2(_2467_),
    .B(_1243_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6855_ (.I(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6856_ (.A1(_2338_),
    .A2(_2467_),
    .B1(_2517_),
    .B2(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6857_ (.A1(_2476_),
    .A2(_2504_),
    .B(_2520_),
    .C(_2293_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6858_ (.A1(_2463_),
    .A2(_2521_),
    .B(_2045_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6859_ (.A1(_1689_),
    .A2(_2359_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6860_ (.A1(\as2650.pc[4] ),
    .A2(_2465_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6861_ (.A1(_1688_),
    .A2(_2523_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _6862_ (.A1(_1592_),
    .A2(_0577_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6863_ (.A1(_2468_),
    .A2(_2470_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6864_ (.A1(_1586_),
    .A2(_0976_),
    .B(_2526_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6865_ (.A1(_2525_),
    .A2(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6866_ (.A1(_2267_),
    .A2(_2528_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6867_ (.A1(_2266_),
    .A2(_2524_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6868_ (.A1(_2474_),
    .A2(_2529_),
    .A3(_2530_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6869_ (.I(_2125_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6870_ (.A1(_2362_),
    .A2(_2531_),
    .B(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6871_ (.I(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6872_ (.I(_1713_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6873_ (.A1(\as2650.stack[1][5] ),
    .A2(_2402_),
    .B1(_2535_),
    .B2(\as2650.stack[0][5] ),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6874_ (.A1(\as2650.stack[3][5] ),
    .A2(_2507_),
    .B1(_2510_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6875_ (.A1(_2506_),
    .A2(_2536_),
    .A3(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6876_ (.A1(\as2650.stack[5][5] ),
    .A2(_1547_),
    .B1(_1651_),
    .B2(\as2650.stack[7][5] ),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6877_ (.A1(\as2650.stack[4][5] ),
    .A2(_2535_),
    .B1(_2400_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6878_ (.A1(_2513_),
    .A2(_2539_),
    .A3(_2540_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6879_ (.A1(_2538_),
    .A2(_2541_),
    .B(_2116_),
    .C(_1264_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6880_ (.A1(_1587_),
    .A2(_2480_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6881_ (.A1(_1593_),
    .A2(_2543_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6882_ (.A1(_1269_),
    .A2(_2056_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6883_ (.A1(_3725_),
    .A2(_2327_),
    .B(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6884_ (.A1(_1520_),
    .A2(_2524_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(_1210_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6886_ (.A1(_2430_),
    .A2(_2528_),
    .B(_2547_),
    .C(_2548_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6887_ (.A1(_2308_),
    .A2(_2544_),
    .B1(_2546_),
    .B2(_1873_),
    .C(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6888_ (.A1(_0495_),
    .A2(_2489_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6889_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_3482_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6890_ (.A1(_0577_),
    .A2(_2552_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6891_ (.A1(_2551_),
    .A2(_2494_),
    .A3(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6892_ (.A1(_2551_),
    .A2(_2494_),
    .B(_2553_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6893_ (.A1(_2059_),
    .A2(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6894_ (.A1(_2554_),
    .A2(_2556_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6895_ (.A1(_1270_),
    .A2(_2493_),
    .B(_2497_),
    .C(_2557_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6896_ (.A1(_2121_),
    .A2(_2550_),
    .B(_2558_),
    .C(_2442_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6897_ (.A1(_1855_),
    .A2(_2524_),
    .B1(_2531_),
    .B2(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6898_ (.A1(_2542_),
    .A2(_2560_),
    .B(_2532_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6899_ (.A1(_2524_),
    .A2(_2534_),
    .B(_2561_),
    .C(_2293_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6900_ (.A1(_2522_),
    .A2(_2562_),
    .B(_2045_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6901_ (.A1(\as2650.pc[6] ),
    .A2(_1688_),
    .A3(_2523_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6902_ (.A1(_1689_),
    .A2(_2523_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6903_ (.A1(_1598_),
    .A2(_2564_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6904_ (.A1(_2563_),
    .A2(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6905_ (.I(_2566_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6906_ (.A1(\as2650.pc[6] ),
    .A2(_0668_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6907_ (.I(_2568_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6908_ (.A1(\as2650.pc[4] ),
    .A2(net9),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6909_ (.A1(_1593_),
    .A2(_1483_),
    .B(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6910_ (.A1(\as2650.pc[5] ),
    .A2(_0577_),
    .B(_2571_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6911_ (.A1(_2468_),
    .A2(_2470_),
    .A3(_2525_),
    .B(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6912_ (.A1(_2569_),
    .A2(_2573_),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6913_ (.A1(_2306_),
    .A2(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6914_ (.A1(_2464_),
    .A2(_2567_),
    .B(_2575_),
    .C(_2475_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6915_ (.A1(_1688_),
    .A2(_1586_),
    .A3(_2480_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6916_ (.A1(_1597_),
    .A2(_2577_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6917_ (.I(_2248_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6918_ (.A1(_2579_),
    .A2(_2566_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6919_ (.I(_2548_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6920_ (.A1(_1521_),
    .A2(_2574_),
    .B(_2580_),
    .C(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6921_ (.I(_2385_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6922_ (.A1(_1424_),
    .A2(_2583_),
    .B1(_1853_),
    .B2(_3605_),
    .C(_2032_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6923_ (.A1(_2250_),
    .A2(_2578_),
    .B1(_2582_),
    .B2(_2584_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6924_ (.I(_2384_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6925_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_3482_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6926_ (.A1(_1454_),
    .A2(_2587_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6927_ (.I(_0668_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6928_ (.A1(_2589_),
    .A2(_2587_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6929_ (.A1(_0578_),
    .A2(_2552_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6930_ (.A1(_2588_),
    .A2(_2590_),
    .B(_2591_),
    .C(_2555_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6931_ (.A1(_2591_),
    .A2(_2555_),
    .B(_2588_),
    .C(_2590_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6932_ (.A1(_2427_),
    .A2(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6933_ (.A1(_2592_),
    .A2(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6934_ (.A1(_1848_),
    .A2(_2586_),
    .B(_2434_),
    .C(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6935_ (.A1(_1945_),
    .A2(_2585_),
    .B(_2596_),
    .C(_2479_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6936_ (.A1(_2478_),
    .A2(_2567_),
    .B1(_2597_),
    .B2(_2503_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6937_ (.I(_2337_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6938_ (.A1(_2599_),
    .A2(_2567_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6939_ (.I(_2284_),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6940_ (.A1(\as2650.stack[0][6] ),
    .A2(_2508_),
    .B1(_2601_),
    .B2(\as2650.stack[2][6] ),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6941_ (.I(_2286_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6942_ (.I(_2283_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6943_ (.A1(\as2650.stack[1][6] ),
    .A2(_2603_),
    .B1(_2604_),
    .B2(\as2650.stack[3][6] ),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6944_ (.A1(_2506_),
    .A2(_2602_),
    .A3(_2605_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6945_ (.A1(\as2650.stack[4][6] ),
    .A2(_2508_),
    .B1(_2601_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6946_ (.A1(\as2650.stack[5][6] ),
    .A2(_2603_),
    .B1(_2604_),
    .B2(\as2650.stack[7][6] ),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6947_ (.A1(_2513_),
    .A2(_2607_),
    .A3(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6948_ (.A1(_2113_),
    .A2(_2606_),
    .A3(_2609_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6949_ (.A1(_2505_),
    .A2(_2567_),
    .B(_2610_),
    .C(_2353_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6950_ (.A1(_2576_),
    .A2(_2598_),
    .B(_2600_),
    .C(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6951_ (.A1(_1691_),
    .A2(_2357_),
    .B(_2461_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6952_ (.A1(_2298_),
    .A2(_2612_),
    .B(_2613_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6953_ (.A1(_1693_),
    .A2(_2563_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6954_ (.I(_2614_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6955_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6956_ (.A1(_1597_),
    .A2(_1454_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6957_ (.A1(_2569_),
    .A2(_2573_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6958_ (.A1(_2617_),
    .A2(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6959_ (.A1(_2616_),
    .A2(_2619_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6960_ (.A1(_2306_),
    .A2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6961_ (.A1(_2464_),
    .A2(_2615_),
    .B(_2621_),
    .C(_2475_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6962_ (.A1(_1598_),
    .A2(_2577_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6963_ (.A1(_1602_),
    .A2(_2623_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6964_ (.A1(_2579_),
    .A2(_2614_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6965_ (.A1(_1521_),
    .A2(_2620_),
    .B(_2625_),
    .C(_2581_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6966_ (.A1(_2216_),
    .A2(_2057_),
    .B1(_1853_),
    .B2(_1850_),
    .C(_2032_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6967_ (.A1(_2250_),
    .A2(_2624_),
    .B1(_2626_),
    .B2(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6968_ (.A1(net3),
    .A2(_3652_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6969_ (.A1(_2588_),
    .A2(_2593_),
    .A3(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6970_ (.A1(_2588_),
    .A2(_2593_),
    .B(_2629_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6971_ (.A1(_2583_),
    .A2(_2631_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6972_ (.A1(_2216_),
    .A2(_2493_),
    .B(_2498_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6973_ (.A1(_2630_),
    .A2(_2632_),
    .B(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6974_ (.A1(_1945_),
    .A2(_2628_),
    .B(_2634_),
    .C(_2246_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6975_ (.A1(_2478_),
    .A2(_2615_),
    .B1(_2635_),
    .B2(_2532_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6976_ (.A1(_2599_),
    .A2(_2615_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6977_ (.A1(\as2650.stack[7][7] ),
    .A2(_2604_),
    .B1(_2601_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6978_ (.A1(\as2650.stack[5][7] ),
    .A2(_2603_),
    .B1(_2535_),
    .B2(\as2650.stack[4][7] ),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6979_ (.A1(_2513_),
    .A2(_2638_),
    .A3(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6980_ (.A1(\as2650.stack[1][7] ),
    .A2(_2603_),
    .B1(_2601_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6981_ (.A1(\as2650.stack[3][7] ),
    .A2(_2604_),
    .B1(_2535_),
    .B2(\as2650.stack[0][7] ),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6982_ (.A1(_2346_),
    .A2(_2641_),
    .A3(_2642_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6983_ (.A1(_2113_),
    .A2(_2640_),
    .A3(_2643_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6984_ (.A1(_2505_),
    .A2(_2615_),
    .B(_2644_),
    .C(_2353_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6985_ (.A1(_2622_),
    .A2(_2636_),
    .B(_2637_),
    .C(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6986_ (.A1(_1694_),
    .A2(_2357_),
    .B(_2461_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6987_ (.A1(_2298_),
    .A2(_2646_),
    .B(_2647_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6988_ (.A1(_1609_),
    .A2(_2359_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6989_ (.A1(\as2650.pc[8] ),
    .A2(_0668_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6990_ (.I(_2649_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6991_ (.A1(_2568_),
    .A2(_2616_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6992_ (.A1(_1693_),
    .A2(_1454_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6993_ (.A1(_2617_),
    .A2(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6994_ (.A1(_2573_),
    .A2(_2651_),
    .B(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6995_ (.A1(_2650_),
    .A2(_2654_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_2650_),
    .A2(_2654_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6997_ (.A1(_2655_),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6998_ (.A1(_1602_),
    .A2(_2563_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6999_ (.A1(_1607_),
    .A2(_2658_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7000_ (.I(_2659_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7001_ (.A1(_2422_),
    .A2(_2657_),
    .B1(_2660_),
    .B2(_2464_),
    .C(_2475_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7002_ (.A1(_0782_),
    .A2(_3652_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7003_ (.A1(_2662_),
    .A2(_2631_),
    .B(_0938_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7004_ (.A1(_2253_),
    .A2(_2663_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7005_ (.A1(_2248_),
    .A2(_2659_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7006_ (.A1(_2380_),
    .A2(_2657_),
    .B(_2665_),
    .C(_1953_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7007_ (.A1(_1412_),
    .A2(_0940_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7008_ (.A1(_1833_),
    .A2(_2059_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7009_ (.A1(_2667_),
    .A2(_2668_),
    .B(_1255_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7010_ (.A1(_1694_),
    .A2(_2623_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7011_ (.A1(_1608_),
    .A2(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7012_ (.A1(_2001_),
    .A2(_2666_),
    .A3(_2669_),
    .B1(_2378_),
    .B2(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7013_ (.A1(_2434_),
    .A2(_2664_),
    .B1(_2672_),
    .B2(_2377_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7014_ (.A1(_2479_),
    .A2(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7015_ (.A1(_2478_),
    .A2(_2660_),
    .B1(_2674_),
    .B2(_2532_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7016_ (.A1(\as2650.stack[7][8] ),
    .A2(_2278_),
    .B1(_2275_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7017_ (.A1(\as2650.stack[5][8] ),
    .A2(_2277_),
    .B1(_2447_),
    .B2(\as2650.stack[4][8] ),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7018_ (.A1(_2444_),
    .A2(_2676_),
    .A3(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_2281_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7020_ (.A1(\as2650.stack[1][8] ),
    .A2(_2277_),
    .B1(_2272_),
    .B2(\as2650.stack[0][8] ),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7021_ (.A1(\as2650.stack[3][8] ),
    .A2(_2278_),
    .B1(_2275_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7022_ (.A1(_2679_),
    .A2(_2680_),
    .A3(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7023_ (.A1(_1218_),
    .A2(_2678_),
    .A3(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7024_ (.A1(_2408_),
    .A2(_2660_),
    .B(_2683_),
    .C(_1243_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7025_ (.I(_2684_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7026_ (.A1(_2599_),
    .A2(_2660_),
    .B(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7027_ (.A1(_2661_),
    .A2(_2675_),
    .B(_2686_),
    .C(_2293_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7028_ (.I(_2044_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7029_ (.A1(_2648_),
    .A2(_2687_),
    .B(_2688_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7030_ (.A1(_1606_),
    .A2(_2658_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7031_ (.A1(_1700_),
    .A2(_2689_),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7032_ (.A1(_1612_),
    .A2(_0669_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7033_ (.A1(_1607_),
    .A2(_1098_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7034_ (.A1(_2692_),
    .A2(_2655_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7035_ (.A1(_2691_),
    .A2(_2693_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7036_ (.A1(_2422_),
    .A2(_2694_),
    .B1(_2690_),
    .B2(_2364_),
    .C(_2474_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7037_ (.A1(_2362_),
    .A2(_2695_),
    .B(_2375_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7038_ (.A1(_2248_),
    .A2(_2690_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7039_ (.A1(_2380_),
    .A2(_2694_),
    .B(_2697_),
    .C(_1953_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7040_ (.A1(_1836_),
    .A2(_2059_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7041_ (.A1(_2330_),
    .A2(_2699_),
    .B(_1255_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7042_ (.A1(_1607_),
    .A2(_1693_),
    .A3(_2623_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7043_ (.A1(_1613_),
    .A2(_2701_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7044_ (.A1(_2001_),
    .A2(_2698_),
    .A3(_2700_),
    .B1(_2702_),
    .B2(_2378_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7045_ (.A1(\as2650.addr_buff[0] ),
    .A2(_2663_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7046_ (.A1(_2314_),
    .A2(_2704_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7047_ (.A1(_2498_),
    .A2(_2705_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7048_ (.A1(_2377_),
    .A2(_2703_),
    .B(_2706_),
    .C(_2442_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7049_ (.A1(\as2650.stack_ptr[2] ),
    .A2(\as2650.stack[3][9] ),
    .B1(_2447_),
    .B2(\as2650.stack[0][9] ),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7050_ (.A1(\as2650.stack[1][9] ),
    .A2(_2451_),
    .B1(_2448_),
    .B2(\as2650.stack[2][9] ),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7051_ (.A1(_2679_),
    .A2(_2708_),
    .A3(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7052_ (.A1(\as2650.stack[5][9] ),
    .A2(_2340_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _7053_ (.A1(\as2650.stack[7][9] ),
    .A2(_2283_),
    .B1(_2284_),
    .B2(\as2650.stack[6][9] ),
    .C1(_1713_),
    .C2(\as2650.stack[4][9] ),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7054_ (.A1(_2444_),
    .A2(_2711_),
    .A3(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7055_ (.A1(_2112_),
    .A2(_2710_),
    .A3(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7056_ (.A1(_2339_),
    .A2(_2690_),
    .B(_2714_),
    .C(_2456_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7057_ (.A1(_2695_),
    .A2(_2707_),
    .B(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7058_ (.A1(_2690_),
    .A2(_2696_),
    .B1(_2716_),
    .B2(_2459_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7059_ (.A1(_2243_),
    .A2(_2717_),
    .B(_2461_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7060_ (.A1(_1614_),
    .A2(_2244_),
    .B(_2718_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7061_ (.A1(_1699_),
    .A2(_1606_),
    .A3(_2658_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7062_ (.A1(_1702_),
    .A2(_2719_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_2305_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7064_ (.A1(\as2650.pc[10] ),
    .A2(_2589_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7065_ (.A1(_1699_),
    .A2(_1606_),
    .B(_2589_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7066_ (.A1(_2655_),
    .A2(_2691_),
    .B(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7067_ (.A1(_2722_),
    .A2(_2724_),
    .Z(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7068_ (.A1(_2721_),
    .A2(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7069_ (.A1(_2364_),
    .A2(_2720_),
    .B(_2726_),
    .C(_2107_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7070_ (.A1(_2247_),
    .A2(_2727_),
    .B(_2126_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7071_ (.A1(_1520_),
    .A2(_2725_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7072_ (.A1(_2430_),
    .A2(_2720_),
    .B(_2729_),
    .C(_1953_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7073_ (.A1(\as2650.addr_buff[2] ),
    .A2(_2385_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7074_ (.A1(_2396_),
    .A2(_2731_),
    .B(_2381_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7075_ (.A1(_1613_),
    .A2(_2701_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7076_ (.A1(_1703_),
    .A2(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7077_ (.A1(_2001_),
    .A2(_2730_),
    .A3(_2732_),
    .B1(_2308_),
    .B2(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7078_ (.A1(_2252_),
    .A2(_2313_),
    .A3(_2383_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7079_ (.A1(_2663_),
    .A2(_2736_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7080_ (.A1(_2314_),
    .A2(_2704_),
    .B(_2383_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7081_ (.A1(_2737_),
    .A2(_2738_),
    .B(_2498_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7082_ (.A1(_2121_),
    .A2(_2735_),
    .B(_2739_),
    .C(_2442_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7083_ (.A1(\as2650.stack[3][10] ),
    .A2(_2445_),
    .B1(_2447_),
    .B2(\as2650.stack[0][10] ),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7084_ (.A1(\as2650.stack[1][10] ),
    .A2(_2451_),
    .B1(_2448_),
    .B2(\as2650.stack[2][10] ),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7085_ (.A1(_2679_),
    .A2(_2741_),
    .A3(_2742_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7086_ (.A1(\as2650.stack[7][10] ),
    .A2(_2445_),
    .B1(_2448_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7087_ (.A1(\as2650.stack[5][10] ),
    .A2(_2451_),
    .B1(_2287_),
    .B2(\as2650.stack[4][10] ),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7088_ (.A1(_2444_),
    .A2(_2744_),
    .A3(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7089_ (.A1(_2112_),
    .A2(_2743_),
    .A3(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7090_ (.A1(_2339_),
    .A2(_2720_),
    .B(_2747_),
    .C(_2456_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7091_ (.A1(_2740_),
    .A2(_2727_),
    .B(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7092_ (.A1(_2720_),
    .A2(_2728_),
    .B1(_2749_),
    .B2(_2459_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7093_ (.I(_0807_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7094_ (.A1(_2243_),
    .A2(_2750_),
    .B(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7095_ (.A1(_1617_),
    .A2(_2244_),
    .B(_2752_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7096_ (.A1(_1616_),
    .A2(_2719_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7097_ (.A1(_1619_),
    .A2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(_2754_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7099_ (.A1(_1702_),
    .A2(_2733_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7100_ (.A1(_1620_),
    .A2(_2756_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7101_ (.I(\as2650.addr_buff[3] ),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7102_ (.A1(_2758_),
    .A2(_2737_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7103_ (.A1(\as2650.addr_buff[3] ),
    .A2(_2663_),
    .A3(_2736_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7104_ (.A1(_2434_),
    .A2(_2759_),
    .A3(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7105_ (.A1(_2247_),
    .A2(_2755_),
    .B1(_2757_),
    .B2(_2251_),
    .C(_2761_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7106_ (.A1(\as2650.pc[11] ),
    .A2(_2589_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7107_ (.A1(\as2650.pc[10] ),
    .A2(_0669_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7108_ (.I(_2722_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7109_ (.A1(_2765_),
    .A2(_2724_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7110_ (.A1(_2764_),
    .A2(_2766_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7111_ (.A1(_2763_),
    .A2(_2767_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7112_ (.A1(_2579_),
    .A2(_2754_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7113_ (.A1(_2579_),
    .A2(_2768_),
    .B(_2769_),
    .C(_2581_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7114_ (.A1(_1841_),
    .A2(_2327_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7115_ (.A1(_2440_),
    .A2(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7116_ (.A1(_1233_),
    .A2(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7117_ (.A1(_2770_),
    .A2(_2773_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7118_ (.A1(_2305_),
    .A2(_2768_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7119_ (.A1(_2363_),
    .A2(_2755_),
    .B(_2775_),
    .C(_2474_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7120_ (.A1(_2246_),
    .A2(_2762_),
    .B1(_2774_),
    .B2(_2090_),
    .C(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7121_ (.A1(\as2650.stack[0][11] ),
    .A2(_2272_),
    .B1(_2343_),
    .B2(\as2650.stack[2][11] ),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7122_ (.A1(\as2650.stack[1][11] ),
    .A2(_2340_),
    .B1(_2278_),
    .B2(\as2650.stack[3][11] ),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7123_ (.A1(_2679_),
    .A2(_2778_),
    .A3(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7124_ (.A1(\as2650.stack[5][11] ),
    .A2(_2340_),
    .B1(_2343_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7125_ (.A1(\as2650.stack[7][11] ),
    .A2(_2342_),
    .B1(_2272_),
    .B2(\as2650.stack[4][11] ),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7126_ (.A1(_2271_),
    .A2(_2781_),
    .A3(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7127_ (.A1(_1218_),
    .A2(_2780_),
    .A3(_2783_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7128_ (.A1(_2408_),
    .A2(_2755_),
    .B(_2784_),
    .C(_2456_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7129_ (.A1(_2375_),
    .A2(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7130_ (.A1(_2503_),
    .A2(_2755_),
    .B1(_2777_),
    .B2(_2786_),
    .C(_2297_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7131_ (.A1(_1621_),
    .A2(_2298_),
    .B(_2787_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7132_ (.A1(_2296_),
    .A2(_2788_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7133_ (.A1(_1619_),
    .A2(_2753_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7134_ (.A1(_1624_),
    .A2(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7135_ (.I(_2790_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7136_ (.A1(_2722_),
    .A2(_2763_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(_2764_),
    .A2(_2723_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7138_ (.A1(\as2650.pc[11] ),
    .A2(_1097_),
    .B(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7139_ (.A1(_2655_),
    .A2(_2691_),
    .A3(_2792_),
    .B(_2794_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7140_ (.A1(\as2650.pc[12] ),
    .A2(_1097_),
    .Z(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7141_ (.A1(_2795_),
    .A2(_2796_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7142_ (.A1(_2721_),
    .A2(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7143_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2385_),
    .B(_2499_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7144_ (.A1(_2365_),
    .A2(_2790_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7145_ (.A1(_1520_),
    .A2(_2797_),
    .B(_1211_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7146_ (.A1(_2548_),
    .A2(_2799_),
    .B1(_2800_),
    .B2(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7147_ (.A1(_2482_),
    .A2(_2760_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7148_ (.A1(_2121_),
    .A2(_2802_),
    .B1(_2803_),
    .B2(_1826_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7149_ (.A1(_1619_),
    .A2(_1702_),
    .A3(_2733_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7150_ (.A1(_1624_),
    .A2(_2805_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7151_ (.A1(_2477_),
    .A2(_2791_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7152_ (.A1(_1446_),
    .A2(_2804_),
    .B1(_2806_),
    .B2(_2251_),
    .C(_2807_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7153_ (.A1(_2266_),
    .A2(_2791_),
    .B1(_2808_),
    .B2(_2246_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7154_ (.A1(_2798_),
    .A2(_2809_),
    .B(_1898_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7155_ (.A1(_1674_),
    .A2(_1711_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7156_ (.A1(_1543_),
    .A2(_1711_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7157_ (.A1(\as2650.stack[5][12] ),
    .A2(_2811_),
    .B1(_2812_),
    .B2(\as2650.stack[7][12] ),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7158_ (.A1(_1543_),
    .A2(_1544_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7159_ (.A1(_1674_),
    .A2(_1544_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7160_ (.A1(\as2650.stack[4][12] ),
    .A2(_2814_),
    .B1(_2815_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7161_ (.A1(_2346_),
    .A2(_2813_),
    .A3(_2816_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7162_ (.A1(\as2650.stack[3][12] ),
    .A2(_2812_),
    .B1(_2815_),
    .B2(\as2650.stack[2][12] ),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7163_ (.A1(\as2650.stack[1][12] ),
    .A2(_2811_),
    .B1(_2814_),
    .B2(\as2650.stack[0][12] ),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7164_ (.A1(_2271_),
    .A2(_2818_),
    .A3(_2819_),
    .B(_2339_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7165_ (.A1(_2505_),
    .A2(_2791_),
    .B1(_2817_),
    .B2(_2820_),
    .C(_2353_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7166_ (.A1(_2297_),
    .A2(_2821_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7167_ (.A1(_2599_),
    .A2(_2791_),
    .B(_2810_),
    .C(_2822_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7168_ (.A1(_1625_),
    .A2(_2357_),
    .B(_2159_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7169_ (.A1(_2823_),
    .A2(_2824_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7170_ (.I(_2384_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7171_ (.I(_1799_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7172_ (.I(_2826_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7173_ (.I(_2827_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7174_ (.A1(_2828_),
    .A2(_3731_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7175_ (.I(_2070_),
    .Z(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7176_ (.A1(_2830_),
    .A2(_3740_),
    .B(_2825_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7177_ (.I(_1328_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7178_ (.I(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7179_ (.A1(_2825_),
    .A2(_3796_),
    .B1(_2829_),
    .B2(_2831_),
    .C(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7180_ (.A1(_0802_),
    .A2(_1229_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7181_ (.I(_2835_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7182_ (.A1(_3767_),
    .A2(_1231_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7183_ (.A1(\as2650.psu[0] ),
    .A2(_2836_),
    .B(_2837_),
    .C(_1445_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7184_ (.I(_1391_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7185_ (.A1(_1379_),
    .A2(_2188_),
    .B1(_3664_),
    .B2(_2839_),
    .C(_1941_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7186_ (.A1(_1453_),
    .A2(_1410_),
    .B1(_2838_),
    .B2(_2840_),
    .C(_1939_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_3553_),
    .A2(_3584_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7188_ (.A1(_1370_),
    .A2(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7189_ (.I(_3556_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7190_ (.A1(_1886_),
    .A2(_2844_),
    .A3(_1330_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7191_ (.A1(_1236_),
    .A2(_1895_),
    .A3(_1344_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7192_ (.A1(_1779_),
    .A2(_0572_),
    .B(_2846_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7193_ (.A1(_3787_),
    .A2(_1266_),
    .A3(_1365_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7194_ (.A1(_1819_),
    .A2(_2304_),
    .A3(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7195_ (.A1(_1327_),
    .A2(_2845_),
    .A3(_2847_),
    .A4(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7196_ (.A1(_3607_),
    .A2(_0973_),
    .B1(_1310_),
    .B2(_1901_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7197_ (.A1(_1808_),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7198_ (.A1(_3537_),
    .A2(_3562_),
    .A3(_1896_),
    .A4(_1797_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7199_ (.A1(_3553_),
    .A2(_3610_),
    .B1(_2852_),
    .B2(_1318_),
    .C(_2853_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7200_ (.A1(_2171_),
    .A2(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7201_ (.A1(_2843_),
    .A2(_2850_),
    .A3(_2855_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7202_ (.I(_2856_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7203_ (.I(_1819_),
    .Z(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7204_ (.I(_2161_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7205_ (.A1(_2858_),
    .A2(_3692_),
    .B1(_2859_),
    .B2(_3784_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7206_ (.A1(_2857_),
    .A2(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7207_ (.I(_2857_),
    .Z(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7208_ (.A1(_2834_),
    .A2(_2841_),
    .A3(_2861_),
    .B1(_2862_),
    .B2(_0865_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7209_ (.A1(_2296_),
    .A2(_2863_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7210_ (.I(_2856_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7211_ (.I(_2864_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7212_ (.I(_1970_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7213_ (.A1(_1331_),
    .A2(_2000_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7214_ (.I(_2867_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7215_ (.I(_2868_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7216_ (.I(_2075_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7217_ (.A1(_2870_),
    .A2(_3900_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7218_ (.I(_2074_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7219_ (.A1(_2828_),
    .A2(_3908_),
    .B(_2871_),
    .C(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7220_ (.A1(_2866_),
    .A2(_3833_),
    .B(_2869_),
    .C(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7221_ (.I(_3675_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7222_ (.I(_1230_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7223_ (.A1(_1292_),
    .A2(_2876_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7224_ (.I(_2835_),
    .Z(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7225_ (.A1(\as2650.psu[1] ),
    .A2(_2878_),
    .B(_3597_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7226_ (.A1(_1395_),
    .A2(_0883_),
    .B1(_2877_),
    .B2(_2879_),
    .C(_3582_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7227_ (.A1(_1400_),
    .A2(_0960_),
    .B(_1940_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7228_ (.A1(_1416_),
    .A2(_2875_),
    .B1(_2880_),
    .B2(_2881_),
    .C(_2373_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7229_ (.A1(_2116_),
    .A2(_3881_),
    .B(_2882_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7230_ (.A1(_2188_),
    .A2(_2162_),
    .B1(_2883_),
    .B2(_1442_),
    .C(_2864_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7231_ (.A1(_2189_),
    .A2(_2865_),
    .B1(_2874_),
    .B2(_2884_),
    .C(_2131_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7232_ (.I(_2857_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7233_ (.I(_2118_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7234_ (.I(_2826_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7235_ (.A1(_2887_),
    .A2(_0321_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7236_ (.A1(_2070_),
    .A2(_0277_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7237_ (.A1(_2886_),
    .A2(_2888_),
    .A3(_2889_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7238_ (.A1(_2872_),
    .A2(_0266_),
    .B(_2868_),
    .C(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7239_ (.A1(_1482_),
    .A2(_2876_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7240_ (.A1(\as2650.overflow ),
    .A2(_1231_),
    .B(_2892_),
    .C(_1444_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7241_ (.A1(_2839_),
    .A2(_2188_),
    .B1(_2197_),
    .B2(_1398_),
    .C(_1940_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7242_ (.A1(_0289_),
    .A2(_2875_),
    .B1(_2893_),
    .B2(_2894_),
    .C(_1938_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7243_ (.A1(_2858_),
    .A2(_0284_),
    .B1(_2859_),
    .B2(_0887_),
    .C(_2895_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7244_ (.A1(_2862_),
    .A2(_2891_),
    .A3(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7245_ (.A1(_2016_),
    .A2(_2885_),
    .B(_2897_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7246_ (.A1(_2296_),
    .A2(_2898_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7247_ (.I(_2044_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7248_ (.A1(_2887_),
    .A2(_0380_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7249_ (.A1(_2887_),
    .A2(_0376_),
    .B(_2900_),
    .C(_1970_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7250_ (.A1(_2872_),
    .A2(_0368_),
    .B(_2868_),
    .C(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7251_ (.A1(_3644_),
    .A2(_2878_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7252_ (.A1(\as2650.psu[3] ),
    .A2(_2836_),
    .B(_2903_),
    .C(_1444_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7253_ (.A1(_2839_),
    .A2(_0887_),
    .B1(_0449_),
    .B2(_1398_),
    .C(_1940_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7254_ (.A1(_1840_),
    .A2(_2875_),
    .B1(_2904_),
    .B2(_2905_),
    .C(_1938_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7255_ (.A1(_2858_),
    .A2(_0384_),
    .B1(_2161_),
    .B2(_2197_),
    .C(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7256_ (.A1(_2857_),
    .A2(_2902_),
    .A3(_2907_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7257_ (.A1(_2020_),
    .A2(_2885_),
    .B(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7258_ (.A1(_2899_),
    .A2(_2909_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7259_ (.A1(_2828_),
    .A2(_0491_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7260_ (.A1(_2830_),
    .A2(_0517_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7261_ (.A1(_2872_),
    .A2(_2910_),
    .A3(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7262_ (.A1(_2866_),
    .A2(_0972_),
    .B(_2869_),
    .C(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7263_ (.I(_2858_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7264_ (.A1(_3650_),
    .A2(_2878_),
    .B(_1392_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7265_ (.A1(\as2650.psu[4] ),
    .A2(_2836_),
    .B(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7266_ (.A1(_0707_),
    .A2(_2197_),
    .B(_2052_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7267_ (.A1(_1379_),
    .A2(_1096_),
    .B1(_2916_),
    .B2(_2917_),
    .C(_1409_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7268_ (.A1(_1423_),
    .A2(_1941_),
    .B(_2918_),
    .C(_1939_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7269_ (.A1(_2914_),
    .A2(_0494_),
    .B1(_2162_),
    .B2(_0561_),
    .C(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7270_ (.A1(_2913_),
    .A2(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7271_ (.A1(_2028_),
    .A2(_2862_),
    .B(_2751_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7272_ (.A1(_2885_),
    .A2(_2921_),
    .B(_2922_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7273_ (.A1(_2830_),
    .A2(_0588_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7274_ (.A1(_2828_),
    .A2(_0559_),
    .B(_2886_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7275_ (.A1(_2825_),
    .A2(_0553_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7276_ (.A1(_2923_),
    .A2(_2924_),
    .B(_2869_),
    .C(_2925_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7277_ (.A1(_1392_),
    .A2(_0449_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7278_ (.A1(_1457_),
    .A2(_2878_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7279_ (.A1(\as2650.psu[5] ),
    .A2(_2836_),
    .B(_2928_),
    .C(_1395_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7280_ (.A1(_2927_),
    .A2(_2929_),
    .B(_1400_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7281_ (.A1(_1400_),
    .A2(_0706_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7282_ (.A1(_1375_),
    .A2(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7283_ (.A1(_1271_),
    .A2(_1375_),
    .B1(_2930_),
    .B2(_2932_),
    .C(_2409_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7284_ (.A1(_2409_),
    .A2(_0576_),
    .B(_2933_),
    .C(_1374_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7285_ (.A1(_0663_),
    .A2(_1364_),
    .B(_2926_),
    .C(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7286_ (.A1(_1017_),
    .A2(_2862_),
    .B(_2751_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7287_ (.A1(_2885_),
    .A2(_2935_),
    .B(_2936_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7288_ (.A1(_2070_),
    .A2(_0679_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7289_ (.A1(_2870_),
    .A2(_0660_),
    .B(_2886_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7290_ (.I(_2867_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7291_ (.A1(_2866_),
    .A2(_1055_),
    .B1(_2937_),
    .B2(_2938_),
    .C(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7292_ (.A1(_1485_),
    .A2(_2876_),
    .B(_2052_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7293_ (.A1(_1388_),
    .A2(_1231_),
    .B(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7294_ (.A1(_1398_),
    .A2(_1101_),
    .B1(_0663_),
    .B2(_1392_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7295_ (.A1(_2942_),
    .A2(_2943_),
    .B(_1409_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7296_ (.A1(_1424_),
    .A2(_1941_),
    .B(_2944_),
    .C(_1939_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7297_ (.A1(_2914_),
    .A2(_0667_),
    .B1(_2859_),
    .B2(_0775_),
    .C(_2945_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7298_ (.A1(_2940_),
    .A2(_2946_),
    .B(_2865_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7299_ (.I(_2044_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7300_ (.A1(_1380_),
    .A2(_2865_),
    .B(_2947_),
    .C(_2948_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7301_ (.A1(_2870_),
    .A2(_0774_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7302_ (.A1(_2830_),
    .A2(_0790_),
    .B(_2886_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7303_ (.A1(_2866_),
    .A2(_1436_),
    .B1(_2949_),
    .B2(_2950_),
    .C(_2939_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7304_ (.A1(\as2650.psl[7] ),
    .A2(_1230_),
    .B(_1377_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7305_ (.A1(_1481_),
    .A2(_2876_),
    .B(_2952_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7306_ (.A1(_1394_),
    .A2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7307_ (.A1(_1399_),
    .A2(_2954_),
    .B(_1409_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7308_ (.A1(_2216_),
    .A2(_2875_),
    .B(_2955_),
    .C(_1938_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7309_ (.A1(_2914_),
    .A2(_0780_),
    .B1(_2859_),
    .B2(_1401_),
    .C(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7310_ (.A1(_2951_),
    .A2(_2957_),
    .B(_2864_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7311_ (.A1(_1114_),
    .A2(_2865_),
    .B(_2958_),
    .C(_2948_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7312_ (.A1(_1628_),
    .A2(_2400_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7313_ (.I(_2959_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7314_ (.I(_2960_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7315_ (.I(_2960_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7316_ (.A1(\as2650.stack[7][0] ),
    .A2(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7317_ (.A1(_1709_),
    .A2(_2961_),
    .B(_2963_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7318_ (.I(_2959_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7319_ (.I0(_1679_),
    .I1(\as2650.stack[7][1] ),
    .S(_2964_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7320_ (.I(_2965_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7321_ (.I0(_1681_),
    .I1(\as2650.stack[7][2] ),
    .S(_2964_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7322_ (.I(_2966_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7323_ (.I(_2960_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7324_ (.A1(\as2650.stack[7][3] ),
    .A2(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7325_ (.A1(_1723_),
    .A2(_2961_),
    .B(_2968_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7326_ (.I(_2960_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7327_ (.I0(_1685_),
    .I1(\as2650.stack[7][4] ),
    .S(_2969_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7328_ (.I(_2970_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7329_ (.A1(\as2650.stack[7][5] ),
    .A2(_2967_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7330_ (.A1(_1594_),
    .A2(_2961_),
    .B(_2971_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7331_ (.A1(\as2650.stack[7][6] ),
    .A2(_2967_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7332_ (.A1(_1599_),
    .A2(_2961_),
    .B(_2972_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7333_ (.A1(\as2650.stack[7][7] ),
    .A2(_2967_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7334_ (.A1(_1603_),
    .A2(_2962_),
    .B(_2973_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7335_ (.I0(_1696_),
    .I1(\as2650.stack[7][8] ),
    .S(_2969_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7336_ (.I(_2974_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7337_ (.A1(\as2650.stack[7][9] ),
    .A2(_2964_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7338_ (.A1(_1732_),
    .A2(_2962_),
    .B(_2975_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7339_ (.A1(\as2650.stack[7][10] ),
    .A2(_2964_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7340_ (.A1(_1734_),
    .A2(_2962_),
    .B(_2976_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7341_ (.I0(_1705_),
    .I1(\as2650.stack[7][11] ),
    .S(_2969_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7342_ (.I(_2977_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7343_ (.I0(_1707_),
    .I1(\as2650.stack[7][12] ),
    .S(_2969_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7344_ (.I(_2978_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7345_ (.A1(_1023_),
    .A2(_3731_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7346_ (.A1(_1413_),
    .A2(_2979_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7347_ (.A1(_3736_),
    .A2(_3734_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7348_ (.A1(_2981_),
    .A2(_3740_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7349_ (.A1(_1413_),
    .A2(_2982_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7350_ (.I(_1802_),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7351_ (.A1(_2870_),
    .A2(_2980_),
    .B1(_2983_),
    .B2(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7352_ (.A1(_1919_),
    .A2(_1794_),
    .A3(_1239_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7353_ (.I(_2986_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7354_ (.I(net28),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7355_ (.A1(_2137_),
    .A2(_2254_),
    .B1(_2987_),
    .B2(_2988_),
    .C(_2832_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7356_ (.A1(_1921_),
    .A2(_2985_),
    .B(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7357_ (.A1(_2053_),
    .A2(_1385_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7358_ (.I(_2991_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7359_ (.A1(_2581_),
    .A2(_2333_),
    .B(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7360_ (.A1(_1352_),
    .A2(_2304_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7361_ (.I(_2994_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7362_ (.A1(_2988_),
    .A2(_2427_),
    .B(_2257_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7363_ (.A1(_2333_),
    .A2(_2254_),
    .B1(_2995_),
    .B2(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7364_ (.A1(_2107_),
    .A2(_1528_),
    .A3(_2997_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7365_ (.A1(_1673_),
    .A2(_2993_),
    .B(_2998_),
    .C(_1433_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7366_ (.A1(_2990_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7367_ (.A1(_1870_),
    .A2(_1364_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7368_ (.I(_3001_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7369_ (.A1(_1194_),
    .A2(_1926_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7370_ (.A1(_3003_),
    .A2(_1930_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7371_ (.A1(_1791_),
    .A2(_1827_),
    .B(_1906_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7372_ (.A1(_3846_),
    .A2(_1968_),
    .A3(_1898_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7373_ (.A1(_3005_),
    .A2(_3006_),
    .B(_1195_),
    .C(_2304_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7374_ (.A1(_1789_),
    .A2(_1504_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7375_ (.A1(_1981_),
    .A2(_3008_),
    .B(_2236_),
    .C(_1822_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7376_ (.A1(_1266_),
    .A2(_1201_),
    .B1(_3003_),
    .B2(_1933_),
    .C(_3009_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7377_ (.A1(_1918_),
    .A2(_1908_),
    .A3(_2225_),
    .A4(_3010_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7378_ (.A1(_1894_),
    .A2(_3007_),
    .A3(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7379_ (.A1(_3004_),
    .A2(_3012_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7380_ (.I(_3013_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7381_ (.A1(_1937_),
    .A2(_3000_),
    .B1(_3002_),
    .B2(_1673_),
    .C(_3014_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7382_ (.A1(_3004_),
    .A2(_3012_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7383_ (.I(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7384_ (.I(_3017_),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7385_ (.A1(_2988_),
    .A2(_3018_),
    .B(_2159_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7386_ (.A1(_3015_),
    .A2(_3019_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7387_ (.I(_3017_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7388_ (.A1(_1990_),
    .A2(_2161_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7389_ (.I(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7390_ (.A1(_1232_),
    .A2(_2305_),
    .B(_2473_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7391_ (.I(_3023_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7392_ (.A1(net52),
    .A2(net28),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7393_ (.A1(_0940_),
    .A2(_3025_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7394_ (.A1(_2315_),
    .A2(_3026_),
    .B(_2994_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7395_ (.A1(_2048_),
    .A2(_2303_),
    .B(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7396_ (.A1(_2992_),
    .A2(_3028_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7397_ (.A1(_1571_),
    .A2(_3024_),
    .B(_3029_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7398_ (.I(_1800_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7399_ (.I(_2844_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7400_ (.A1(_0315_),
    .A2(_1913_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7401_ (.I(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7402_ (.A1(_3665_),
    .A2(_3739_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _7403_ (.A1(_1458_),
    .A2(_3893_),
    .A3(_3905_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7404_ (.A1(_3035_),
    .A2(_3036_),
    .B(_2981_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7405_ (.A1(_3035_),
    .A2(_3036_),
    .B(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7406_ (.A1(_1415_),
    .A2(_3032_),
    .B(_3034_),
    .C(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7407_ (.I(_0314_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7408_ (.A1(_3665_),
    .A2(_3730_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _7409_ (.A1(_1459_),
    .A2(_3893_),
    .A3(_3897_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7410_ (.A1(_3041_),
    .A2(_3042_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7411_ (.I(_0313_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7412_ (.A1(_3041_),
    .A2(_3042_),
    .B(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7413_ (.A1(_1415_),
    .A2(_3040_),
    .B1(_3043_),
    .B2(_3045_),
    .C(_2069_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7414_ (.A1(_1919_),
    .A2(_1890_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7415_ (.A1(_3039_),
    .A2(_3046_),
    .B(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7416_ (.I(_1796_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7417_ (.A1(_3031_),
    .A2(_3025_),
    .B(_3048_),
    .C(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7418_ (.I(_2078_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7419_ (.A1(_1535_),
    .A2(net5),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7420_ (.A1(_3052_),
    .A2(_2302_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7421_ (.A1(_3051_),
    .A2(_3053_),
    .B(_2833_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7422_ (.A1(_1374_),
    .A2(_3030_),
    .B1(_3050_),
    .B2(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7423_ (.I(_1990_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7424_ (.A1(_1572_),
    .A2(_3022_),
    .B1(_3055_),
    .B2(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7425_ (.I(_3017_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7426_ (.A1(net52),
    .A2(_3058_),
    .B(_2751_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7427_ (.A1(_3020_),
    .A2(_3057_),
    .B(_3059_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7428_ (.I(net30),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7429_ (.I(_3013_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7430_ (.A1(_1990_),
    .A2(_2832_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7431_ (.A1(net52),
    .A2(_2988_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7432_ (.A1(_3060_),
    .A2(_3063_),
    .Z(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7433_ (.A1(_2987_),
    .A2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7434_ (.I(_2981_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _7435_ (.A1(_1459_),
    .A2(_3906_),
    .A3(_3907_),
    .B1(_3035_),
    .B2(_3036_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7436_ (.A1(_0270_),
    .A2(_0276_),
    .B(_0287_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7437_ (.A1(_1417_),
    .A2(_0277_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7438_ (.A1(_3068_),
    .A2(_3069_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7439_ (.I(_2844_),
    .Z(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7440_ (.A1(_3067_),
    .A2(_3070_),
    .B(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7441_ (.A1(_3067_),
    .A2(_3070_),
    .B(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7442_ (.A1(_1418_),
    .A2(_3066_),
    .B(_2984_),
    .C(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _7443_ (.A1(_1459_),
    .A2(_3898_),
    .A3(_3899_),
    .B1(_3041_),
    .B2(_3042_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7444_ (.A1(_0317_),
    .A2(_0320_),
    .B(_0288_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7445_ (.A1(_1417_),
    .A2(_0321_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7446_ (.A1(_3076_),
    .A2(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7447_ (.A1(_3075_),
    .A2(_3078_),
    .B(_3044_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7448_ (.A1(_3075_),
    .A2(_3078_),
    .B(_3079_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7449_ (.A1(_1418_),
    .A2(_1024_),
    .B(_2827_),
    .C(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7450_ (.A1(_3074_),
    .A2(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7451_ (.A1(_3052_),
    .A2(_2302_),
    .B(_2366_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7452_ (.A1(_2368_),
    .A2(_3083_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7453_ (.I(_2078_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7454_ (.A1(_1795_),
    .A2(_3082_),
    .B1(_3084_),
    .B2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7455_ (.A1(_3065_),
    .A2(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7456_ (.A1(_3062_),
    .A2(_3087_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7457_ (.A1(_2074_),
    .A2(_3064_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7458_ (.A1(_2386_),
    .A2(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7459_ (.A1(_2991_),
    .A2(_2994_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7460_ (.I(_3091_),
    .Z(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7461_ (.A1(_3090_),
    .A2(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7462_ (.I(_3023_),
    .Z(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7463_ (.A1(_1577_),
    .A2(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7464_ (.A1(_2372_),
    .A2(_3093_),
    .A3(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7465_ (.A1(_1578_),
    .A2(_3002_),
    .B1(_3096_),
    .B2(_2127_),
    .C(_3014_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7466_ (.A1(_3060_),
    .A2(_3061_),
    .B1(_3088_),
    .B2(_3097_),
    .C(_2131_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7467_ (.A1(net30),
    .A2(net52),
    .A3(net28),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7468_ (.A1(net31),
    .A2(_3098_),
    .Z(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7469_ (.A1(_2327_),
    .A2(_3099_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7470_ (.A1(_1421_),
    .A2(_2057_),
    .B(_2995_),
    .C(_3100_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7471_ (.A1(_2048_),
    .A2(_2421_),
    .B(_3101_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7472_ (.A1(_1683_),
    .A2(_1233_),
    .A3(_2721_),
    .B1(_3102_),
    .B2(_2035_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7473_ (.A1(_0287_),
    .A2(_0317_),
    .A3(_0320_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7474_ (.A1(_3075_),
    .A2(_3076_),
    .B(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7475_ (.A1(_0388_),
    .A2(_0380_),
    .A3(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7476_ (.A1(_3044_),
    .A2(_3106_),
    .B(_2075_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7477_ (.A1(_1421_),
    .A2(_3040_),
    .B(_3107_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7478_ (.A1(_0287_),
    .A2(_0270_),
    .A3(_0276_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7479_ (.A1(_3067_),
    .A2(_3068_),
    .B(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7480_ (.A1(_1420_),
    .A2(_0376_),
    .A3(_3110_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7481_ (.A1(_1472_),
    .A2(_3066_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7482_ (.A1(_3066_),
    .A2(_3111_),
    .B(_3112_),
    .C(_3034_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7483_ (.I(_3047_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7484_ (.A1(_3108_),
    .A2(_3113_),
    .B(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7485_ (.I(_2077_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7486_ (.A1(_2986_),
    .A2(_3099_),
    .B(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7487_ (.A1(_2368_),
    .A2(_3083_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7488_ (.A1(_2419_),
    .A2(_3118_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7489_ (.A1(_2418_),
    .A2(_3119_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7490_ (.A1(_2099_),
    .A2(_3120_),
    .B(_2867_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7491_ (.A1(_3115_),
    .A2(_3117_),
    .B(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7492_ (.A1(_1582_),
    .A2(_1812_),
    .B1(_2914_),
    .B2(_3103_),
    .C(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7493_ (.A1(_1683_),
    .A2(_3022_),
    .B1(_3123_),
    .B2(_3056_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7494_ (.I(_0807_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7495_ (.A1(net31),
    .A2(_3058_),
    .B(_3125_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7496_ (.A1(_3020_),
    .A2(_3124_),
    .B(_3126_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7497_ (.I(_2468_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7498_ (.A1(\as2650.pc[3] ),
    .A2(_0386_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7499_ (.A1(_2416_),
    .A2(_3119_),
    .B(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7500_ (.A1(_3127_),
    .A2(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7501_ (.A1(_0387_),
    .A2(_0379_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7502_ (.A1(_0387_),
    .A2(_0379_),
    .B1(_3075_),
    .B2(_3076_),
    .C(_3104_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7503_ (.A1(_1479_),
    .A2(_0491_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7504_ (.A1(_3131_),
    .A2(_3132_),
    .B(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7505_ (.A1(_3131_),
    .A2(_3133_),
    .A3(_3132_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7506_ (.A1(_3044_),
    .A2(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7507_ (.A1(_1480_),
    .A2(_3040_),
    .B1(_3134_),
    .B2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7508_ (.A1(_0275_),
    .A2(_0371_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7509_ (.A1(_0372_),
    .A2(_0373_),
    .B(_3138_),
    .C(_0374_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7510_ (.A1(_0387_),
    .A2(_3139_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7511_ (.A1(_0386_),
    .A2(_3139_),
    .B1(_3067_),
    .B2(_3068_),
    .C(_3109_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7512_ (.A1(_3140_),
    .A2(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7513_ (.A1(_1479_),
    .A2(_0517_),
    .A3(_3142_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7514_ (.A1(_3071_),
    .A2(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7515_ (.A1(_1480_),
    .A2(_3032_),
    .B(_3033_),
    .C(_3144_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7516_ (.A1(_2827_),
    .A2(_3137_),
    .B(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7517_ (.I(net32),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7518_ (.I(net31),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7519_ (.A1(_3148_),
    .A2(_3098_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7520_ (.A1(_3147_),
    .A2(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7521_ (.A1(_1921_),
    .A2(_3146_),
    .B1(_3150_),
    .B2(_1800_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7522_ (.A1(_3051_),
    .A2(_3130_),
    .B(_3151_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7523_ (.A1(_2427_),
    .A2(_3150_),
    .B(_2485_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7524_ (.A1(_2245_),
    .A2(_2471_),
    .B1(_2995_),
    .B2(_3153_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7525_ (.A1(_2373_),
    .A2(_1528_),
    .A3(_3154_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7526_ (.A1(_1587_),
    .A2(_2993_),
    .B(_3155_),
    .C(_1433_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7527_ (.A1(_2833_),
    .A2(_3152_),
    .B(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7528_ (.A1(_1588_),
    .A2(_3002_),
    .B1(_3157_),
    .B2(_1937_),
    .C(_3014_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7529_ (.I(_1430_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7530_ (.A1(_3147_),
    .A2(_3058_),
    .B(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7531_ (.A1(_3158_),
    .A2(_3160_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7532_ (.A1(_3147_),
    .A2(_3149_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7533_ (.A1(net51),
    .A2(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7534_ (.A1(_1477_),
    .A2(_0516_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7535_ (.A1(_1478_),
    .A2(_0516_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7536_ (.A1(_3140_),
    .A2(_3163_),
    .A3(_3141_),
    .B(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7537_ (.A1(_1846_),
    .A2(_0559_),
    .A3(_3165_),
    .Z(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7538_ (.A1(_1269_),
    .A2(_3071_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7539_ (.A1(_3032_),
    .A2(_3166_),
    .B(_3167_),
    .C(_2984_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7540_ (.A1(_0580_),
    .A2(_0588_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7541_ (.A1(_1478_),
    .A2(_0490_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7542_ (.A1(_1478_),
    .A2(_0490_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7543_ (.A1(_3131_),
    .A2(_3170_),
    .A3(_3132_),
    .B(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7544_ (.A1(_3169_),
    .A2(_3172_),
    .B(_0314_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7545_ (.A1(_3169_),
    .A2(_3172_),
    .B(_3173_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7546_ (.A1(_1846_),
    .A2(_1024_),
    .B(_2827_),
    .C(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7547_ (.A1(_3168_),
    .A2(_3175_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7548_ (.A1(_3114_),
    .A2(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7549_ (.A1(_3031_),
    .A2(_3162_),
    .B(_3177_),
    .C(_3049_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7550_ (.A1(_3127_),
    .A2(_3129_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7551_ (.A1(_2570_),
    .A2(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7552_ (.A1(_2525_),
    .A2(_3180_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7553_ (.A1(_3051_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7554_ (.A1(_3062_),
    .A2(_3178_),
    .A3(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7555_ (.I(_3091_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7556_ (.A1(_2074_),
    .A2(_3162_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7557_ (.A1(_2545_),
    .A2(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7558_ (.A1(_1689_),
    .A2(_3024_),
    .B1(_3184_),
    .B2(_3186_),
    .C(_2338_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7559_ (.A1(_1593_),
    .A2(_3001_),
    .B1(_3187_),
    .B2(_2529_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7560_ (.A1(_3183_),
    .A2(_3188_),
    .B(_3061_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7561_ (.A1(net51),
    .A2(_3058_),
    .B(_3159_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7562_ (.A1(_3189_),
    .A2(_3190_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7563_ (.A1(net51),
    .A2(_3147_),
    .A3(_3149_),
    .ZN(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7564_ (.A1(net34),
    .A2(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7565_ (.A1(_1424_),
    .A2(_2583_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7566_ (.A1(_2586_),
    .A2(_3192_),
    .B(_3193_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7567_ (.A1(_1691_),
    .A2(_3024_),
    .B1(_3184_),
    .B2(_3194_),
    .C(_1319_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7568_ (.A1(_2525_),
    .A2(_3179_),
    .B(_2572_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7569_ (.A1(_2569_),
    .A2(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7570_ (.A1(_1456_),
    .A2(_0678_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7571_ (.A1(_0579_),
    .A2(_0587_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7572_ (.A1(_0579_),
    .A2(_0587_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7573_ (.A1(_3199_),
    .A2(_3172_),
    .B(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7574_ (.A1(_3198_),
    .A2(_3201_),
    .B(_0314_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7575_ (.A1(_3198_),
    .A2(_3201_),
    .B(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7576_ (.A1(_1848_),
    .A2(_1023_),
    .B(_2826_),
    .C(_3203_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7577_ (.A1(_1455_),
    .A2(_0659_),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7578_ (.A1(_0578_),
    .A2(_0558_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7579_ (.A1(_0578_),
    .A2(_0558_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7580_ (.A1(_3165_),
    .A2(_3206_),
    .B(_3207_),
    .ZN(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7581_ (.A1(_3205_),
    .A2(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7582_ (.A1(_2981_),
    .A2(_3209_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7583_ (.A1(_1456_),
    .A2(_3066_),
    .B(_1802_),
    .C(_3210_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7584_ (.A1(_3204_),
    .A2(_3211_),
    .B(_2167_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7585_ (.A1(_2986_),
    .A2(_3192_),
    .B(_3212_),
    .C(_3116_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7586_ (.A1(_3085_),
    .A2(_3197_),
    .B(_3213_),
    .C(_2833_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7587_ (.A1(_2575_),
    .A2(_3195_),
    .B(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7588_ (.A1(_1691_),
    .A2(_3022_),
    .B1(_3215_),
    .B2(_3056_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7589_ (.I(_3016_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7590_ (.A1(net34),
    .A2(_3217_),
    .B(_3125_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7591_ (.A1(_3020_),
    .A2(_3216_),
    .B(_3218_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7592_ (.I(net35),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7593_ (.A1(net34),
    .A2(net51),
    .A3(net32),
    .A4(_3149_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7594_ (.A1(_3219_),
    .A2(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7595_ (.A1(_0670_),
    .A2(_0679_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7596_ (.A1(_3198_),
    .A2(_3201_),
    .B(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7597_ (.A1(_1981_),
    .A2(_0790_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7598_ (.A1(_3223_),
    .A2(_3224_),
    .B(_1023_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7599_ (.A1(_3223_),
    .A2(_3224_),
    .B(_3225_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7600_ (.A1(_1449_),
    .A2(_3040_),
    .B(_2069_),
    .C(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7601_ (.A1(_1097_),
    .A2(_0660_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7602_ (.A1(_3205_),
    .A2(_3208_),
    .B(_3228_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7603_ (.A1(_1115_),
    .A2(_0774_),
    .A3(_3229_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7604_ (.A1(_3071_),
    .A2(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7605_ (.A1(_1449_),
    .A2(_3032_),
    .B(_3034_),
    .C(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7606_ (.A1(_3227_),
    .A2(_3232_),
    .B(_3047_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7607_ (.A1(_3031_),
    .A2(_3221_),
    .B(_3233_),
    .C(_3049_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7608_ (.A1(_2569_),
    .A2(_3196_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7609_ (.A1(_2617_),
    .A2(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7610_ (.A1(_2616_),
    .A2(_3236_),
    .B(_2099_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7611_ (.A1(_2616_),
    .A2(_3236_),
    .B(_3237_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7612_ (.A1(_3062_),
    .A2(_3234_),
    .A3(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7613_ (.I0(_1449_),
    .I1(_3221_),
    .S(_2118_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7614_ (.A1(_1694_),
    .A2(_3094_),
    .B1(_3092_),
    .B2(_3240_),
    .C(_2337_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7615_ (.A1(_1602_),
    .A2(_3001_),
    .B1(_3241_),
    .B2(_2621_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7616_ (.A1(_3239_),
    .A2(_3242_),
    .B(_3014_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7617_ (.A1(_3219_),
    .A2(_3061_),
    .B(_3243_),
    .C(_2948_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7618_ (.A1(_2651_),
    .A2(_3196_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7619_ (.A1(_2617_),
    .A2(_2652_),
    .A3(_3244_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7620_ (.A1(_2649_),
    .A2(_3245_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7621_ (.A1(_2649_),
    .A2(_3245_),
    .B(_3085_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7622_ (.A1(_1115_),
    .A2(_0789_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7623_ (.A1(_3198_),
    .A2(_3201_),
    .B(_3248_),
    .C(_3222_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7624_ (.A1(_1981_),
    .A2(_0789_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7625_ (.A1(_0313_),
    .A2(_3250_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7626_ (.A1(_1833_),
    .A2(_3249_),
    .A3(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7627_ (.A1(_3249_),
    .A2(_3251_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7628_ (.A1(_2253_),
    .A2(_3253_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7629_ (.A1(_3252_),
    .A2(_3254_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7630_ (.A1(_0782_),
    .A2(_0773_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7631_ (.A1(_3205_),
    .A2(_3208_),
    .B(_3256_),
    .C(_3228_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7632_ (.A1(_1115_),
    .A2(_0773_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7633_ (.A1(_2844_),
    .A2(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7634_ (.A1(\as2650.addr_buff[0] ),
    .A2(_3257_),
    .A3(_3259_),
    .ZN(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7635_ (.A1(_3257_),
    .A2(_3259_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7636_ (.A1(_2253_),
    .A2(_3261_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7637_ (.A1(_3260_),
    .A2(_3262_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7638_ (.A1(_2887_),
    .A2(_3255_),
    .B1(_3263_),
    .B2(_2984_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7639_ (.A1(_3219_),
    .A2(_3220_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7640_ (.A1(net50),
    .A2(_3265_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7641_ (.I(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7642_ (.A1(_2986_),
    .A2(_3267_),
    .B(_3116_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7643_ (.A1(_2167_),
    .A2(_3264_),
    .B(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7644_ (.A1(_3246_),
    .A2(_3247_),
    .B(_2939_),
    .C(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7645_ (.A1(_2721_),
    .A2(_2657_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7646_ (.A1(_2586_),
    .A2(_3267_),
    .B(_3091_),
    .C(_2668_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7647_ (.A1(_1608_),
    .A2(_2993_),
    .B(_3271_),
    .C(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7648_ (.A1(_2503_),
    .A2(_3273_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7649_ (.A1(_1609_),
    .A2(_3021_),
    .B1(_3270_),
    .B2(_1991_),
    .C(_3274_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7650_ (.A1(net50),
    .A2(_3217_),
    .B(_3125_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7651_ (.A1(_3020_),
    .A2(_3275_),
    .B(_3276_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7652_ (.A1(_1699_),
    .A2(_0670_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7653_ (.A1(_1608_),
    .A2(_1387_),
    .B(_3246_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7654_ (.A1(_3277_),
    .A2(_3278_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7655_ (.A1(net50),
    .A2(_3265_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7656_ (.A1(net37),
    .A2(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7657_ (.A1(_2314_),
    .A2(_3260_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7658_ (.A1(_3034_),
    .A2(_3282_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7659_ (.A1(_1836_),
    .A2(_3252_),
    .B(_2075_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7660_ (.A1(_1836_),
    .A2(_3252_),
    .B(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7661_ (.A1(_3283_),
    .A2(_3285_),
    .B(_3047_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7662_ (.A1(_3031_),
    .A2(_3281_),
    .B(_3286_),
    .C(_2099_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7663_ (.A1(_3049_),
    .A2(_3279_),
    .B(_3287_),
    .C(_2939_),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7664_ (.A1(_2493_),
    .A2(_3281_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7665_ (.A1(_2699_),
    .A2(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7666_ (.A1(_1700_),
    .A2(_3094_),
    .B1(_3092_),
    .B2(_3290_),
    .C(_2337_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7667_ (.A1(_2422_),
    .A2(_2694_),
    .B(_3291_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7668_ (.A1(_1700_),
    .A2(_3021_),
    .B1(_3288_),
    .B2(_1991_),
    .C(_3292_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7669_ (.A1(net37),
    .A2(_3217_),
    .B(_3125_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7670_ (.A1(_3018_),
    .A2(_3293_),
    .B(_3294_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7671_ (.A1(net37),
    .A2(net50),
    .A3(_3265_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7672_ (.A1(net38),
    .A2(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7673_ (.A1(_2586_),
    .A2(_3296_),
    .B(_2731_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7674_ (.A1(_1703_),
    .A2(_3024_),
    .B1(_3184_),
    .B2(_3297_),
    .C(_1319_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7675_ (.A1(_3257_),
    .A2(_3259_),
    .B(_2826_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7676_ (.A1(_1913_),
    .A2(_2736_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7677_ (.A1(_3249_),
    .A2(_3251_),
    .B(_2069_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7678_ (.A1(_1833_),
    .A2(\as2650.addr_buff[1] ),
    .B(_1801_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7679_ (.A1(_1914_),
    .A2(_3299_),
    .B(_3301_),
    .C(_3302_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7680_ (.A1(_3299_),
    .A2(_3300_),
    .A3(_3301_),
    .B1(_3303_),
    .B2(\as2650.addr_buff[2] ),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7681_ (.A1(_3114_),
    .A2(_3304_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7682_ (.A1(_2987_),
    .A2(_3296_),
    .B(_3116_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7683_ (.I(_2723_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7684_ (.A1(_3277_),
    .A2(_3246_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7685_ (.A1(_2765_),
    .A2(_3307_),
    .A3(_3308_),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7686_ (.A1(_3307_),
    .A2(_3308_),
    .B(_2765_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7687_ (.A1(_3309_),
    .A2(_3310_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7688_ (.A1(_3305_),
    .A2(_3306_),
    .B1(_3311_),
    .B2(_2137_),
    .C(_2832_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7689_ (.A1(_2726_),
    .A2(_3298_),
    .B(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7690_ (.A1(_1703_),
    .A2(_3022_),
    .B1(_3313_),
    .B2(_3056_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7691_ (.A1(net38),
    .A2(_3217_),
    .B(_1883_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7692_ (.A1(_3018_),
    .A2(_3314_),
    .B(_3315_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7693_ (.I(net38),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7694_ (.A1(_3316_),
    .A2(_3295_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7695_ (.A1(net39),
    .A2(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7696_ (.A1(_2987_),
    .A2(_3318_),
    .B(_2137_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7697_ (.A1(_1801_),
    .A2(_2736_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7698_ (.A1(_1914_),
    .A2(_3299_),
    .B(_3301_),
    .C(_3320_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7699_ (.A1(_2758_),
    .A2(_3299_),
    .A3(_3300_),
    .A4(_3301_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7700_ (.A1(_1841_),
    .A2(_3321_),
    .B(_3322_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7701_ (.A1(_3114_),
    .A2(_3323_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7702_ (.A1(_2764_),
    .A2(_3310_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7703_ (.A1(_2763_),
    .A2(_3325_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7704_ (.A1(_3319_),
    .A2(_3324_),
    .B1(_3326_),
    .B2(_3085_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7705_ (.A1(_2869_),
    .A2(_3327_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7706_ (.A1(_2825_),
    .A2(_3318_),
    .B(_2771_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7707_ (.A1(_3184_),
    .A2(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7708_ (.A1(_1620_),
    .A2(_1322_),
    .A3(_2479_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7709_ (.A1(_1620_),
    .A2(_2992_),
    .B(_2338_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7710_ (.A1(_2775_),
    .A2(_3330_),
    .A3(_3331_),
    .A4(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7711_ (.A1(_1621_),
    .A2(_3021_),
    .B1(_3328_),
    .B2(_1991_),
    .C(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7712_ (.A1(net39),
    .A2(_3017_),
    .B(_1883_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7713_ (.A1(_3018_),
    .A2(_3334_),
    .B(_3335_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7714_ (.I(net40),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7715_ (.A1(net39),
    .A2(_3317_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7716_ (.A1(net40),
    .A2(_3337_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7717_ (.A1(_2758_),
    .A2(_1914_),
    .B(_1844_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7718_ (.A1(_1844_),
    .A2(_3322_),
    .B1(_3321_),
    .B2(_3339_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7719_ (.A1(_1801_),
    .A2(_3338_),
    .B(_3340_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7720_ (.A1(_2765_),
    .A2(_2763_),
    .A3(_3308_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7721_ (.A1(_2794_),
    .A2(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7722_ (.A1(_2796_),
    .A2(_3343_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7723_ (.A1(_1870_),
    .A2(_2868_),
    .ZN(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7724_ (.A1(_2167_),
    .A2(_3338_),
    .B1(_3344_),
    .B2(_3051_),
    .C(_3345_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7725_ (.A1(_1921_),
    .A2(_3341_),
    .B(_3346_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7726_ (.A1(_1844_),
    .A2(_2057_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7727_ (.A1(_2583_),
    .A2(_3338_),
    .B(_3348_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7728_ (.A1(_1624_),
    .A2(_3094_),
    .B1(_3092_),
    .B2(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7729_ (.A1(_2798_),
    .A2(_3350_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7730_ (.A1(_1625_),
    .A2(_3002_),
    .B1(_3351_),
    .B2(_2459_),
    .C(_3013_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7731_ (.A1(_3336_),
    .A2(_3061_),
    .B1(_3347_),
    .B2(_3352_),
    .C(_1986_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7732_ (.A1(_1158_),
    .A2(_1159_),
    .A3(_0412_),
    .A4(_0801_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7733_ (.I(_3353_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7734_ (.A1(_0807_),
    .A2(_3353_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7735_ (.I(_3355_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7736_ (.A1(_3745_),
    .A2(_3356_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7737_ (.A1(_3798_),
    .A2(_3354_),
    .B(_3357_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7738_ (.A1(_3839_),
    .A2(_3356_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7739_ (.A1(_3913_),
    .A2(_3354_),
    .B(_3358_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7740_ (.A1(_3866_),
    .A2(_3356_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7741_ (.A1(_0335_),
    .A2(_3354_),
    .B(_3359_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7742_ (.A1(_0299_),
    .A2(_3356_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7743_ (.A1(_0430_),
    .A2(_3354_),
    .B(_3360_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7744_ (.I(_3353_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7745_ (.I(_3355_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7746_ (.A1(_0394_),
    .A2(_3362_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7747_ (.A1(_0521_),
    .A2(_3361_),
    .B(_3363_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7748_ (.A1(_0500_),
    .A2(_3362_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7749_ (.A1(_0616_),
    .A2(_3361_),
    .B(_3364_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7750_ (.A1(\as2650.r123[0][6] ),
    .A2(_3362_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7751_ (.A1(_0713_),
    .A2(_3361_),
    .B(_3365_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7752_ (.A1(\as2650.r123[0][7] ),
    .A2(_3362_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7753_ (.A1(_0795_),
    .A2(_3361_),
    .B(_3366_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7754_ (.A1(_2992_),
    .A2(_2226_),
    .A3(_2995_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7755_ (.A1(_2430_),
    .A2(_2473_),
    .A3(_2548_),
    .A4(_1818_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7756_ (.A1(_1214_),
    .A2(_1560_),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7757_ (.A1(_2473_),
    .A2(_3369_),
    .B(_2098_),
    .C(_1326_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7758_ (.A1(_3368_),
    .A2(_2323_),
    .A3(_2228_),
    .A4(_3370_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7759_ (.A1(_3612_),
    .A2(_1356_),
    .A3(_1506_),
    .A4(_1976_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7760_ (.A1(_2230_),
    .A2(_3367_),
    .A3(_3371_),
    .A4(_3372_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7761_ (.A1(_1711_),
    .A2(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7762_ (.A1(_2899_),
    .A2(_3374_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7763_ (.I(_3373_),
    .Z(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7764_ (.A1(_2812_),
    .A2(_2815_),
    .B(_2409_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7765_ (.A1(_2108_),
    .A2(_2507_),
    .A3(_2510_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7766_ (.A1(_3376_),
    .A2(_3377_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7767_ (.A1(_1674_),
    .A2(_3375_),
    .B(_1883_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7768_ (.A1(_3375_),
    .A2(_3378_),
    .B(_3379_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7769_ (.A1(_2506_),
    .A2(_3376_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7770_ (.A1(\as2650.stack_ptr[2] ),
    .A2(_3375_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7771_ (.A1(_3375_),
    .A2(_3380_),
    .B(_3381_),
    .C(_2948_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7772_ (.A1(_0860_),
    .A2(_1871_),
    .A3(_1512_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7773_ (.A1(_2108_),
    .A2(_3382_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7774_ (.A1(_1840_),
    .A2(_3382_),
    .B(_3383_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7775_ (.A1(_1434_),
    .A2(_3382_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7776_ (.A1(_1843_),
    .A2(_3382_),
    .B(_3384_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7777_ (.I(_1258_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7778_ (.A1(_3385_),
    .A2(_1268_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7779_ (.A1(_1444_),
    .A2(_2033_),
    .A3(_3386_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7780_ (.A1(_2927_),
    .A2(_2931_),
    .A3(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7781_ (.A1(_1270_),
    .A2(_1299_),
    .A3(_2221_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7782_ (.A1(_3855_),
    .A2(_3639_),
    .B(_3644_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7783_ (.A1(_1995_),
    .A2(_1343_),
    .A3(_2174_),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7784_ (.A1(_1507_),
    .A2(_1208_),
    .B(_2222_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7785_ (.A1(_3772_),
    .A2(_1780_),
    .B(_1252_),
    .C(_1226_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7786_ (.A1(_1354_),
    .A2(_1860_),
    .A3(_3392_),
    .A4(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7787_ (.A1(_1357_),
    .A2(_3394_),
    .ZN(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7788_ (.A1(_3390_),
    .A2(_3391_),
    .A3(_3395_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7789_ (.A1(_2068_),
    .A2(_3388_),
    .B(_3389_),
    .C(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7790_ (.A1(_1434_),
    .A2(_0972_),
    .B(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7791_ (.A1(_3396_),
    .A2(_3389_),
    .B(_1457_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7792_ (.A1(_1884_),
    .A2(_3398_),
    .A3(_3399_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7793_ (.I(_3400_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7794_ (.A1(_1996_),
    .A2(_1401_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7795_ (.A1(_0737_),
    .A2(_1996_),
    .B(_3401_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7796_ (.A1(_0456_),
    .A2(_0457_),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7797_ (.A1(_0698_),
    .A2(_3852_),
    .B(_3762_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7798_ (.A1(_3805_),
    .A2(_3831_),
    .B(_3404_),
    .C(_3795_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7799_ (.A1(_1284_),
    .A2(_3832_),
    .B(_3405_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7800_ (.A1(_0265_),
    .A2(_0353_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7801_ (.A1(_0265_),
    .A2(_0353_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7802_ (.A1(_0363_),
    .A2(_0936_),
    .B1(_3406_),
    .B2(_3407_),
    .C(_3408_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7803_ (.A1(_0363_),
    .A2(_0936_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7804_ (.A1(_3403_),
    .A2(_0465_),
    .B(_3409_),
    .C(_3410_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7805_ (.A1(_3403_),
    .A2(_0465_),
    .B1(_0552_),
    .B2(_0694_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7806_ (.A1(_0552_),
    .A2(_0694_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7807_ (.A1(_0711_),
    .A2(_0723_),
    .B1(_3411_),
    .B2(_3412_),
    .C(_3413_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7808_ (.A1(_1055_),
    .A2(_0723_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7809_ (.A1(_1154_),
    .A2(_3402_),
    .B(_3414_),
    .C(_3415_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7810_ (.A1(_1154_),
    .A2(_3402_),
    .B(_1374_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7811_ (.A1(_1414_),
    .A2(_2015_),
    .A3(_2221_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7812_ (.A1(_3396_),
    .A2(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7813_ (.A1(_3385_),
    .A2(_2008_),
    .B(_2007_),
    .C(_1445_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7814_ (.A1(_1379_),
    .A2(_0883_),
    .B1(_1401_),
    .B2(_2839_),
    .C(_1319_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7815_ (.A1(_3420_),
    .A2(_3421_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7816_ (.A1(_3419_),
    .A2(_3422_),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7817_ (.A1(_3416_),
    .A2(_3417_),
    .B(_3423_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7818_ (.A1(_3767_),
    .A2(_3419_),
    .B(_3159_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7819_ (.A1(_3424_),
    .A2(_3425_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7820_ (.A1(_1436_),
    .A2(_3402_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7821_ (.A1(_1442_),
    .A2(_0731_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7822_ (.A1(_1419_),
    .A2(_2015_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7823_ (.A1(_2107_),
    .A2(_1445_),
    .B(_3391_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7824_ (.A1(_2068_),
    .A2(_3428_),
    .B(_3394_),
    .C(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7825_ (.A1(_3385_),
    .A2(_2017_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7826_ (.A1(_2068_),
    .A2(_2018_),
    .A3(_3431_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7827_ (.A1(_3430_),
    .A2(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7828_ (.A1(_3426_),
    .A2(_3427_),
    .B(_3433_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7829_ (.A1(\as2650.overflow ),
    .A2(_3430_),
    .B(_3159_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7830_ (.A1(_3434_),
    .A2(_3435_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7831_ (.A1(_0803_),
    .A2(_1465_),
    .B1(_1256_),
    .B2(_1507_),
    .C(_1200_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7832_ (.A1(_2006_),
    .A2(_1348_),
    .B(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7833_ (.A1(_1204_),
    .A2(_1254_),
    .A3(_1873_),
    .A4(_3437_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7834_ (.A1(_1843_),
    .A2(_2023_),
    .B(_3438_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7835_ (.A1(_2035_),
    .A2(_3385_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7836_ (.A1(_2028_),
    .A2(_2036_),
    .B(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7837_ (.A1(_3484_),
    .A2(_3439_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7838_ (.A1(_3439_),
    .A2(_3441_),
    .B(_3442_),
    .C(_2132_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7839_ (.A1(_2022_),
    .A2(_2214_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7840_ (.A1(_3443_),
    .A2(_3438_),
    .B(\as2650.psl[3] ),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7841_ (.A1(_2020_),
    .A2(_1967_),
    .B1(_3440_),
    .B2(_2022_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7842_ (.A1(_3438_),
    .A2(_3445_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7843_ (.A1(_3444_),
    .A2(_3446_),
    .B(_2688_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7844_ (.A1(_1460_),
    .A2(_2023_),
    .B(_3438_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7845_ (.A1(_0908_),
    .A2(_2036_),
    .B(_3440_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7846_ (.A1(_1292_),
    .A2(_3447_),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7847_ (.A1(_3447_),
    .A2(_3448_),
    .B(_3449_),
    .C(_2132_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7848_ (.I(_2035_),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7849_ (.A1(_0803_),
    .A2(_1208_),
    .B(_1877_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7850_ (.A1(_1217_),
    .A2(_1226_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7851_ (.A1(_3536_),
    .A2(_1872_),
    .A3(_3451_),
    .A4(_3452_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7852_ (.A1(_1202_),
    .A2(_1866_),
    .A3(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7853_ (.I(_3454_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7854_ (.I(_3455_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7855_ (.A1(_1425_),
    .A2(_3450_),
    .B(_3456_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7856_ (.I(_1274_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7857_ (.A1(_2023_),
    .A2(_3458_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7858_ (.A1(_0662_),
    .A2(_1529_),
    .B1(_3459_),
    .B2(_1848_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7859_ (.I(_3454_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7860_ (.A1(_1485_),
    .A2(_3457_),
    .B1(_3460_),
    .B2(_3461_),
    .C(_1986_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7861_ (.A1(_1423_),
    .A2(_3450_),
    .B(_3456_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7862_ (.A1(\as2650.psu[4] ),
    .A2(_3462_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7863_ (.A1(_2030_),
    .A2(_3461_),
    .A3(_3459_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7864_ (.A1(_3463_),
    .A2(_3464_),
    .B(_2688_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7865_ (.A1(_2022_),
    .A2(_3450_),
    .B(_3455_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7866_ (.A1(_3458_),
    .A2(_2024_),
    .B(_2021_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7867_ (.A1(\as2650.psu[3] ),
    .A2(_3465_),
    .B1(_3466_),
    .B2(_3461_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7868_ (.A1(_2899_),
    .A2(_3467_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7869_ (.A1(_1419_),
    .A2(_2011_),
    .B(_3455_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7870_ (.A1(_1967_),
    .A2(_3458_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7871_ (.A1(_2016_),
    .A2(_2214_),
    .B(_3469_),
    .C(_3468_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7872_ (.A1(_1482_),
    .A2(_3468_),
    .B(_3470_),
    .C(_2132_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7873_ (.A1(_1416_),
    .A2(_3450_),
    .B(_3456_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7874_ (.A1(\as2650.psu[1] ),
    .A2(_3471_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7875_ (.A1(_2013_),
    .A2(_3456_),
    .A3(_3459_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7876_ (.A1(_3472_),
    .A2(_3473_),
    .B(_2688_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7877_ (.A1(_1414_),
    .A2(_2214_),
    .B(_3455_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7878_ (.A1(_3458_),
    .A2(_2008_),
    .B(_2007_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7879_ (.A1(\as2650.psu[0] ),
    .A2(_3474_),
    .B1(_3475_),
    .B2(_3461_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7880_ (.A1(_2899_),
    .A2(_3476_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7881_ (.D(_0000_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7882_ (.D(_0001_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7883_ (.D(_0002_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7884_ (.D(_0003_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7885_ (.D(_0004_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7886_ (.D(_0005_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7887_ (.D(_0006_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7888_ (.D(_0007_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7889_ (.D(_0008_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7890_ (.D(_0009_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7891_ (.D(_0010_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7892_ (.D(_0011_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7893_ (.D(_0012_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7894_ (.D(_0013_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7895_ (.D(_0014_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7896_ (.D(_0015_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7897_ (.D(_0016_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7898_ (.D(_0017_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7899_ (.D(_0018_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7900_ (.D(_0019_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7901_ (.D(_0020_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7902_ (.D(_0021_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7903_ (.D(_0022_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7904_ (.D(_0023_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7905_ (.D(_0024_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7906_ (.D(_0025_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7907_ (.D(_0026_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7908_ (.D(_0027_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7909_ (.D(_0028_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7910_ (.D(_0029_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7911_ (.D(_0030_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7912_ (.D(_0031_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7913_ (.D(_0032_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7914_ (.D(_0033_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7915_ (.D(_0034_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7916_ (.D(_0035_),
    .CLK(clknet_opt_2_0_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7917_ (.D(_0036_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7918_ (.D(_0037_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7919_ (.D(_0038_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7920_ (.D(_0039_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7921_ (.D(_0040_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7922_ (.D(_0041_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7923_ (.D(_0042_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7924_ (.D(_0043_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7925_ (.D(_0044_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7926_ (.D(_0045_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7927_ (.D(_0046_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7928_ (.D(_0047_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7929_ (.D(_0048_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7930_ (.D(_0049_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7931_ (.D(_0050_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7932_ (.D(_0051_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7933_ (.D(_0052_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7934_ (.D(_0053_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7935_ (.D(_0054_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7936_ (.D(_0055_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7937_ (.D(_0056_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7938_ (.D(_0057_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7939_ (.D(_0058_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7940_ (.D(_0059_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7941_ (.D(_0060_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7942_ (.D(_0061_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7943_ (.D(_0062_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7944_ (.D(_0063_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7945_ (.D(_0064_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7946_ (.D(_0065_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7947_ (.D(_0066_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7948_ (.D(_0067_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7949_ (.D(_0068_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7950_ (.D(_0069_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7951_ (.D(_0070_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7952_ (.D(_0071_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7953_ (.D(_0072_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7954_ (.D(_0073_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7955_ (.D(_0074_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7956_ (.D(_0075_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7957_ (.D(_0076_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7958_ (.D(_0077_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7959_ (.D(_0078_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7960_ (.D(_0079_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7961_ (.D(_0080_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7962_ (.D(_0081_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7963_ (.D(_0082_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7964_ (.D(_0083_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7965_ (.D(_0084_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7966_ (.D(_0085_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7967_ (.D(_0086_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7968_ (.D(_0087_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7969_ (.D(_0088_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7970_ (.D(_0089_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7971_ (.D(_0090_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7972_ (.D(_0091_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7973_ (.D(_0092_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7974_ (.D(_0093_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7975_ (.D(_0094_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7976_ (.D(_0095_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7977_ (.D(_0096_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7978_ (.D(_0097_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7979_ (.D(_0098_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7980_ (.D(_0099_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7981_ (.D(_0100_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7982_ (.D(_0101_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7983_ (.D(_0102_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7984_ (.D(_0103_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7985_ (.D(_0104_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7986_ (.D(_0105_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7987_ (.D(_0106_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7988_ (.D(_0107_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7989_ (.D(_0108_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7990_ (.D(_0109_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7991_ (.D(_0110_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7992_ (.D(_0111_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7993_ (.D(_0112_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7994_ (.D(_0113_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7995_ (.D(_0114_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7996_ (.D(_0115_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7997_ (.D(_0116_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7998_ (.D(_0117_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7999_ (.D(_0118_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8000_ (.D(_0119_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8001_ (.D(_0120_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8002_ (.D(_0121_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8003_ (.D(_0122_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8004_ (.D(_0123_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8005_ (.D(_0124_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8006_ (.D(_0125_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8007_ (.D(_0126_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8008_ (.D(_0127_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8009_ (.D(_0128_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8010_ (.D(_0129_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8011_ (.D(_0130_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8012_ (.D(_0131_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8013_ (.D(_0132_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8014_ (.D(_0133_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8015_ (.D(_0134_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8016_ (.D(_0135_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8017_ (.D(_0136_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8018_ (.D(_0137_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8019_ (.D(_0138_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8020_ (.D(_0139_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8021_ (.D(_0140_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8022_ (.D(_0141_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8023_ (.D(_0142_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8024_ (.D(_0143_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8025_ (.D(_0144_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8026_ (.D(_0145_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8027_ (.D(_0146_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8028_ (.D(_0147_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8029_ (.D(_0148_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8030_ (.D(_0149_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8031_ (.D(_0150_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8032_ (.D(_0151_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8033_ (.D(_0152_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8034_ (.D(_0153_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8035_ (.D(_0154_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8036_ (.D(_0155_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8037_ (.D(_0156_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8038_ (.D(_0157_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8039_ (.D(_0158_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8040_ (.D(_0159_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8041_ (.D(_0160_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8042_ (.D(_0161_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8043_ (.D(_0162_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8044_ (.D(_0163_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8045_ (.D(_0164_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8046_ (.D(_0165_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8047_ (.D(_0166_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8048_ (.D(_0167_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8049_ (.D(_0168_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8050_ (.D(_0169_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8051_ (.D(_0170_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8052_ (.D(_0171_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8053_ (.D(_0172_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8054_ (.D(_0173_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8055_ (.D(_0174_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8056_ (.D(_0175_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8057_ (.D(_0176_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8058_ (.D(_0177_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8059_ (.D(_0178_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8060_ (.D(_0179_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8061_ (.D(_0180_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8062_ (.D(_0181_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8063_ (.D(_0182_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8064_ (.D(_0183_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8065_ (.D(_0184_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8066_ (.D(_0185_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8067_ (.D(_0186_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8068_ (.D(_0187_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8069_ (.D(_0188_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8070_ (.D(_0189_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8071_ (.D(_0190_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8072_ (.D(_0191_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8073_ (.D(_0192_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8074_ (.D(_0193_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8075_ (.D(_0194_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8076_ (.D(_0195_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8077_ (.D(_0196_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8078_ (.D(_0197_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8079_ (.D(_0198_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8080_ (.D(_0199_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8081_ (.D(_0200_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8082_ (.D(_0201_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8083_ (.D(_0202_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8084_ (.D(_0203_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8085_ (.D(_0204_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8086_ (.D(_0205_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8087_ (.D(_0206_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8088_ (.D(_0207_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8089_ (.D(_0208_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8090_ (.D(_0209_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8091_ (.D(_0210_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8092_ (.D(_0211_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8093_ (.D(_0212_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8094_ (.D(_0213_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8095_ (.D(_0214_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8096_ (.D(_0215_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8097_ (.D(_0216_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8098_ (.D(_0217_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8099_ (.D(_0218_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8100_ (.D(_0219_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8101_ (.D(_0220_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8102_ (.D(_0221_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8103_ (.D(_0222_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8104_ (.D(_0223_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8105_ (.D(_0224_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8106_ (.D(_0225_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8107_ (.D(_0226_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8108_ (.D(_0227_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8109_ (.D(_0228_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8110_ (.D(_0229_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8111_ (.D(_0230_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8112_ (.D(_0231_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8113_ (.D(_0232_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8114_ (.D(_0233_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8115_ (.D(_0234_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8116_ (.D(_0235_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8117_ (.D(_0236_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8118_ (.D(_0237_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8119_ (.D(_0238_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8120_ (.D(_0239_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8121_ (.D(_0240_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8122_ (.D(_0241_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8123_ (.D(_0242_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8124_ (.D(_0243_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8125_ (.D(_0244_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8126_ (.D(_0245_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8127_ (.D(_0246_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8128_ (.D(_0247_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8129_ (.D(_0248_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8130_ (.D(_0249_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8131_ (.D(_0250_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8132_ (.D(_0251_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8133_ (.D(_0252_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8134_ (.D(_0253_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8135_ (.D(_0254_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8136_ (.D(_0255_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8137_ (.D(_0256_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8138_ (.D(_0257_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8139_ (.D(_0258_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8140_ (.D(_0259_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8141_ (.D(_0260_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_88 (.Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8183_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8184_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8185_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8186_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8187_ (.I(net47),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8188_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8189_ (.I(net47),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[5]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[6]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(io_in[7]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[8]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(io_in[9]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net49),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net13),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net36),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net33),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net29),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_opt_1_1_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_1_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_opt_1_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__D (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__D (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__D (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__D (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__D (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__D (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__D (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__D (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__D (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__D (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__D (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__D (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__D (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__D (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__D (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__D (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__D (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__D (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__D (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__D (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__B2 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__B3 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__C (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__B (.I(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I0 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__C (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__C (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A3 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A3 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__B1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__B1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__A1 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__A1 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__B2 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__I (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__B1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__B2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__B (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__B1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__B1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I0 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A4 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A3 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__C (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__B (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__B (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A3 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A3 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A4 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__B2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__B2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__C (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__S (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__C (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I0 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__S (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A3 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__C (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__B (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__B2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__B2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__B2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__B2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__I (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__I (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__B2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__I (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__B1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I0 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__S (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__B1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__I (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__B1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A4 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__B (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__B (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__B1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A3 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__C (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__B (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A3 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__B1 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A4 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__C (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7805__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7804__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A3 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A3 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__B1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I0 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__B1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A3 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__I (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__B (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__I1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__C (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__B (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__B1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__B1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__B2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__C (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__B (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__B1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A2 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__I (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A3 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A3 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A3 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__B (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A3 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__B1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__B1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__B1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A3 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__B (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__B (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__B (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__B (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__C (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__I (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__C1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__C (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__B (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7751__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A3 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__B (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A3 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__B1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__B2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A3 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A2 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__B (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__B (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A3 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A4 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__B (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__B (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__B (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__S (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__C (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__I (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__C (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__C (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__B (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__B (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__B (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__B (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__B (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__C (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__I (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__C (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A3 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__B (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__B (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__B (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__B2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__B (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__B (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A3 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__C (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__B (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__B (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__B (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__B2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__B (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__B (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__B (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__C (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__B (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A4 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A4 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__I (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__B (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__I (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__C (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__I (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A3 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I0 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I0 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__I (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__I (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__I (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__B (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__B2 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A3 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__B (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I0 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I0 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A2 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I0 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I0 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A2 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A3 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__C1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__C2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__C (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__I0 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I0 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__B (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__I (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__B (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__S (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__S (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__S (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__S (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__I (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__I (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__B (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A3 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__C (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__B (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__I (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__I (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__B (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__B (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A3 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__B (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A1 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A3 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__C (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__I (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A3 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__C (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A3 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A3 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__C (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__B (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A3 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A2 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__B (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__B1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A3 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__B (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__B (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__B1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__B (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A4 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__I (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__C (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__C (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__B (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__C2 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__B (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__B (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__B (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__B (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__I (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__C (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__C (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__C (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__B1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A3 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A3 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__B1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__B2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__B1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__B (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__B2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__C (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__C (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__C (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A4 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A3 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__B2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__B (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__B2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__B1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A3 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A4 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A3 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A4 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A3 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__C (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A3 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A3 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__I (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A2 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__C (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__C (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__C (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A3 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__B (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__C (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__B (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__I (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__C (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__B2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__B2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__B (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__B (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__B (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__C (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__B (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__B1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__B2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__I (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A3 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A1 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__I (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A1 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__I (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A3 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__I (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A4 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__B2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A3 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A4 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7529__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__B (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__B (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__B (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__B (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__C (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__C (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__C (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__I (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__I (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__C (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__C (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__C (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A3 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__B2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__B2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__C (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__C (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__C (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__C (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A1 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__I (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__I (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I0 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__B (.I(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__A1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__B1 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__B (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__B2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A3 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__I (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7541__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__I (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__I (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__B1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__B2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__I (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__B1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__B2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A4 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__I (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__B2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A4 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__B (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__I0 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__B2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__I (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__B (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A3 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__I (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A3 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A3 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__B2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__B (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__B (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A3 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__B1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__C (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A3 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__I (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__B1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__B (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__B2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A3 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__C (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__I (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__B (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__I (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__I (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__I0 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__I0 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__I0 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I0 (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__S (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__S (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__B (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__I (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I0 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__I0 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__I0 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__I0 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__S (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__S (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__S (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__S (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__I (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__I (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__I (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__I (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__I (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__I (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__I (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I0 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__I0 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__I0 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__I0 (.I(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__I (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__S (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__S (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__B1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A3 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__S (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__S (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__S (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__S (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__S (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__S (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__B2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__B2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__S (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__S (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__S (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__S (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__S (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__I0 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__I0 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I0 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__I1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__S (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__S (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__S (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__S (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__I1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__S (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__S (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__S (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__S (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__I1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__I0 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I0 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__I0 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__C1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__B1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__C1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__B1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__B1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A2 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__S (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__S (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__S (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__S (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__S (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__S (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__I (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__I (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__S (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__S (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__S (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__S (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__S (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__S (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__I (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__S (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__S (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__S (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__C (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__I (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A3 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__I (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__I (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A3 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A4 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__I (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A3 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__I (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A1 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A3 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A3 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A4 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A3 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A4 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A3 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__B2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__I (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7583__B (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__I (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A4 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A3 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__B (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__I (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__B (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__I (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__I (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__I (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A4 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__I (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__B (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__C (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__C (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__B (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A3 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__C (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A3 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A4 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__I (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__I (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__I (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__S (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__B (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__B2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__I1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__B1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__B1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__B1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__I (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B1 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__I (.I(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__B2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A3 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A3 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A3 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A3 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A3 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A2 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__B (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__B (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__C (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__I (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__C (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B1 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__C (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A3 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A3 (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__I (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__I (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A2 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__I (.I(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A3 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__B2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__B2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__B (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__I (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__B2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__B (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__B (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A3 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__B (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__B (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__B (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__C (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__I (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A3 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__B (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A2 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A3 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A3 (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A2 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A3 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A3 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__B2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A3 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__B (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A3 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__B2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__B (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__B (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__B (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__B (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__B (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__C (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A2 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__I (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__B (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A3 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__I (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__C (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A4 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__B (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A2 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A3 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__B2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__C (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__C (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__C (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__I (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__C (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__I (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__I (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__C (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__I (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__C (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__B (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__B1 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__C (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__C (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__C (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__C (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__B (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__B1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__I (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__I (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__C (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__B2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__B (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A4 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__C (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__B (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A3 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__C (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__C (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__I (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__I (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__I (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__B2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__B2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__I (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B1 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__S (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__I (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__I (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__S (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__S (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__A1 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__B2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__I (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__B (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__B (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__I0 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__I (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__I0 (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__A1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__B (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__B2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A1 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__I0 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__S (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__S (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__S (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I0 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__C (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__C (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A2 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__I0 (.I(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__I (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__B2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__I (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I0 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I0 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__B (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__B (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__B (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__B (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__B (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__I (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__C (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A3 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__B (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__B (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__B (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__B (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__I (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A2 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__I (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__I (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__C (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__C (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__B (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__B (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A2 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__B (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__B (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__C (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__C (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__B (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__B (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__I (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__B (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A3 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__I (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__I (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__B (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A4 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A3 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A3 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A4 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A1 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A3 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__B2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A2 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__C (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__B (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A1 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__C (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A3 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__I (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__A1 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A3 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__B (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__C (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__S (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__B (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__I (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__I (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__B2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__B2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__C (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__B1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__B2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__C (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__C (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__C (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__C (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__C (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__C (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__C (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__B1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__B (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__B2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A3 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__B (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__B (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__B1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__I (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__B1 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A4 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__B (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__B (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__B1 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A3 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__I (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__I (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__A2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__B2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__B1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__I0 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__I0 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A3 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A3 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A4 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A3 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__C (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A3 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A3 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A3 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A4 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__B (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A3 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A4 (.I(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A4 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__I (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__I (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__I (.I(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__I (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__C (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__I (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A2 (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__I (.I(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__B2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__C (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A2 (.I(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__I (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__B (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__C (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__B (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A2 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__B1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__B1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__B1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__B1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__B1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A2 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__B1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__B1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__B1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__I (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__B1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__I (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__B1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__I (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__B1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__B1 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A2 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__C (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__C (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__C (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__C (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__B1 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__C (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A2 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__I (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__I (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__B2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__B1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A2 (.I(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A2 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__C (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__I (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__C (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__B (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__I (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__C (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__C (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__C (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__B (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__C (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__B (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__B1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__B1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__B1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__B1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__B (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__C (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__C (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__C (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__B2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A2 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A2 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__I (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__B (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A3 (.I(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__B (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__C (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__C (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__C (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A1 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A2 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__B (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__B (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__B (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__B2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__B2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__B1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__B (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__B2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__C (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__C (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__B (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A3 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__C (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__C (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__B (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__B (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A2 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__B1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__B1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__B1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__B (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__C (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__B (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__A2 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__B1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__B2 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A2 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__B1 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__B (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__B (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__C (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__C (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__C (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__C (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A2 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__A1 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__B1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__B1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__B1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__B1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__B1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__B1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__B1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__B1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__B (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__C (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__C (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__C (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__C (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__B2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__B2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__B2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__I (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A2 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__A2 (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__B (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__I (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__C (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__C (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__I (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A3 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__C (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A3 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__B (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__I (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__B1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__B2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__B2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__A2 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A3 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__B1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__B1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A2 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A3 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__B1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__A2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A3 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__B2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A2 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__B1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A3 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__I (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6886__C (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A2 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__B (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__B2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6900__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__B (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__A2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__C (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__C (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__C (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A1 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__B2 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A1 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A2 (.I(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__B (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__C (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__B (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__B1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__B1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__B1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__B1 (.I(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__B1 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__B1 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A3 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__B (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A2 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__B2 (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__B (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__B2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__B (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__B (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__A2 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__B (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__I (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A1 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A3 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A2 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__B1 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__C (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A3 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__B2 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__B1 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__B (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__B (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__B (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__B (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__B (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__B1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__A1 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A2 (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A3 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__B1 (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__B (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__B (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__A2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A1 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__A3 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__B (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__B (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A2 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A3 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__B2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A3 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__B (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A2 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__I (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__B1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A3 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__C (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__B (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__B1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__B (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__I (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A2 (.I(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A1 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B1 (.I(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__B1 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B1 (.I(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__B2 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__B (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__B (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__B (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7173__I (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A1 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__C (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__B (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__C (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__I (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__I (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__B2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__B2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__A2 (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A1 (.I(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__I (.I(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__I (.I(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A2 (.I(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A2 (.I(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__B (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A3 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A2 (.I(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__B (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__C (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I (.I(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A2 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__B (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__B (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A2 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__B (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__B (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__B (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__B (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__B (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__C (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__A2 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A2 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A2 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__B2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__B (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__B (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__B (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__C (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__A3 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__C (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__A2 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__B1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A1 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__B1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A1 (.I(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__C (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__B (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__B (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__C (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__C (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__B (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__C (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__C (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__B (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__C (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A2 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__C (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__C (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__C (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__C (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__B (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__I (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__I (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__I (.I(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__A2 (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__S (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__S (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__S (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__S (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__S (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__S (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__I (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__B (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__B2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__C (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__B (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__B2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__A1 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__I (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__B1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A1 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__B2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A1 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__I (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A1 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__B (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A3 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__B1 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__B (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__B1 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__I (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__B1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A4 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__C (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__I (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__I (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__I (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7692__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A2 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7651__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A2 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__I (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__I (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__I (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A1 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__B (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__I (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__B (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__C (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__B (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__C (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__B1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__A1 (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__B (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__B (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__B2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__B (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__B (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__I (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__B (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__B (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__C (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__C (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__C (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A2 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__B1 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__B (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A1 (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A2 (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__B (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__B2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__B (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__B2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__A2 (.I(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A1 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__B (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__I (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__I (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__B1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__B1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__B1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A2 (.I(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__B2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A2 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7469__A2 (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A3 (.I(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__C (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__B (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__A2 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7681__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__B (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__B (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__B (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__C (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__B (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__C (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__B (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__B (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__B (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__B (.I(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A2 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__B1 (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__B (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__B (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__B (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__B (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__B (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__B2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__A2 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__A2 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__B2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__B (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__B (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__B (.I(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A3 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__B2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__B (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__C (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__C (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__B (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__B (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__B2 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__B2 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__A1 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7688__B1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__B (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__A2 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7704__B1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__B1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A2 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A2 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__B1 (.I(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__C (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__B2 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__B2 (.I(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A2 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A4 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A1 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A2 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__B (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__B (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A3 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__B (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A2 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__C (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7809__B (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A2 (.I(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A2 (.I(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__B (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__B (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A1 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A2 (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__B (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A2 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__I (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__I (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A3 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A3 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__B1 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__B2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__B2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__B2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A2 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A2 (.I(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__S0 (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__S (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__I (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__I (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__S0 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__S0 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__S (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A1 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I (.I(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A3 (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A4 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__I (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__B2 (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__S1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__S1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__B (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__S1 (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__B (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__I (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__I (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__S (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A1 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__I (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A3 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__I (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__I (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A3 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__C (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__I (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__I (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A2 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__I (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A3 (.I(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__C (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__I (.I(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__I (.I(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__I (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__I (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A1 (.I(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__I (.I(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__B2 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__B2 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__I (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__B2 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__B2 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A3 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__B2 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A4 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A1 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__S1 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__I (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A1 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__A2 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A3 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__I (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A2 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__I (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__I (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__C (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__C (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__I (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A3 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__A3 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__I (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A1 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A3 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A3 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__I (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A4 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A3 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A3 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A3 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__I (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A3 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A3 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A1 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__I (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__I (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__I (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__I (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A3 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A3 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A1 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A3 (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__C (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A3 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A2 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__I (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A3 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A3 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A3 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__A1 (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__I (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__I (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__I (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__B (.I(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__I (.I(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A3 (.I(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A2 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__I (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A2 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__B2 (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__B2 (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__B2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A2 (.I(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A2 (.I(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__I (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A2 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A4 (.I(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__A3 (.I(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__S1 (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__S1 (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__I (.I(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A2 (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__I (.I(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__A3 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__I (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__I (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A1 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__B (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__I (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__I (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A3 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__I (.I(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__C (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__I (.I(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__A1 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A2 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__A4 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__I (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__I (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A2 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__B (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A1 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A1 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__I (.I(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A1 (.I(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__B2 (.I(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__I (.I(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__I (.I(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__B (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__B2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__B (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__B1 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A2 (.I(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__A1 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__I (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__I (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__I (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__I (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__I (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__I (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__I (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__I (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__I (.I(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__B (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__C (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__I (.I(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__B2 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__I (.I(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__B1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__B1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A2 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A2 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__B2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__B2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__I (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A1 (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__B1 (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__I (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__B2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__I (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__I (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A1 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__I (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A3 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__I (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__I (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__C (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A1 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__C (.I(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__I (.I(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__B2 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A2 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__A1 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A2 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A1 (.I(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A2 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__B1 (.I(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__B2 (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__B2 (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A3 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A3 (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__I (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__C (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A3 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__B (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__I (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__I (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__I (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__C (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__I (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__I (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__B (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__B (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__B (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__C (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__B2 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__B1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__I (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7818__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A2 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__C (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__I (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A2 (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__B (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A1 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__B2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A1 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A4 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__I (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__B (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A1 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__B2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__B2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__B2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__B2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__I1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A1 (.I(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__A1 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A4 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__I (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__C (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__I (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A4 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__B1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__B (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__I (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__B (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__B (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__B2 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__B (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__I (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A2 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__B1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A4 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__I (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__A1 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__B1 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A4 (.I(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__B (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__C (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__I (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A1 (.I(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__I (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__I (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__I (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__B (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__B (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__B (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__B (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__B (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A2 (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__I (.I(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__C (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__I (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B2 (.I(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__B2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__C1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__A1 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I0 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__B1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__C2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__I (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__I (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__I (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__I (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A2 (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__A2 (.I(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A1 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__I (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__B (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__B2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__A2 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__I (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__B (.I(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__C2 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__B2 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__B (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__B1 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__B (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__I (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__B (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__B (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__I1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__C (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__C (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__B (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A4 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__A2 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A3 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__B (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__C (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__C (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__C (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__B2 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__I (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__C (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__I (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__I (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A3 (.I(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__C (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__I (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__I (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__B2 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__I (.I(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__B (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__B (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__S0 (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__I (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__B2 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__B2 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I (.I(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A4 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__A1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I0 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I0 (.I(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__I0 (.I(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I2 (.I(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I0 (.I(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I2 (.I(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__I0 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I2 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__I0 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I2 (.I(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I0 (.I(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I2 (.I(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__I (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__I (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I1 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__I1 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I1 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__I1 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__I1 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I3 (.I(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__I3 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__I1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I3 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I1 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I3 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__I1 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I3 (.I(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__I1 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I3 (.I(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I1 (.I(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I3 (.I(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I1 (.I(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A1 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I0 (.I(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__I0 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I0 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I0 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I0 (.I(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B2 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B2 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__B2 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__B2 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__B2 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__B2 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__C2 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__B2 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__B2 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__B2 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__B2 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__B2 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__I1 (.I(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__B2 (.I(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__B2 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A1 (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A1 (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A1 (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A3 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A3 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7669__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7715__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__I1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__CLK (.I(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__CLK (.I(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__CLK (.I(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__CLK (.I(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__CLK (.I(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__CLK (.I(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_1_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_opt_1_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__CLK (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net88;
 assign io_oeb[13] = net93;
 assign io_oeb[14] = net53;
 assign io_oeb[15] = net54;
 assign io_oeb[16] = net55;
 assign io_oeb[17] = net56;
 assign io_oeb[18] = net57;
 assign io_oeb[19] = net58;
 assign io_oeb[1] = net89;
 assign io_oeb[20] = net59;
 assign io_oeb[21] = net60;
 assign io_oeb[22] = net61;
 assign io_oeb[23] = net62;
 assign io_oeb[24] = net63;
 assign io_oeb[25] = net64;
 assign io_oeb[26] = net65;
 assign io_oeb[27] = net66;
 assign io_oeb[28] = net67;
 assign io_oeb[29] = net68;
 assign io_oeb[2] = net90;
 assign io_oeb[30] = net69;
 assign io_oeb[31] = net70;
 assign io_oeb[32] = net71;
 assign io_oeb[33] = net72;
 assign io_oeb[34] = net73;
 assign io_oeb[35] = net74;
 assign io_oeb[36] = net75;
 assign io_oeb[37] = net76;
 assign io_oeb[3] = net91;
 assign io_oeb[4] = net92;
 assign io_out[0] = net77;
 assign io_out[13] = net82;
 assign io_out[1] = net78;
 assign io_out[2] = net79;
 assign io_out[33] = net83;
 assign io_out[34] = net84;
 assign io_out[35] = net85;
 assign io_out[36] = net86;
 assign io_out[37] = net87;
 assign io_out[3] = net80;
 assign io_out[4] = net81;
endmodule

