magic
tech gf180mcuD
magscale 1 10
timestamp 1698834931
<< nwell >>
rect 1258 155584 218710 156448
rect 1258 154016 218710 154880
rect 1258 152448 218710 153312
rect 1258 150880 218710 151744
rect 1258 149312 218710 150176
rect 1258 147744 218710 148608
rect 1258 146176 218710 147040
rect 1258 144608 218710 145472
rect 1258 143040 218710 143904
rect 1258 141472 218710 142336
rect 1258 139904 218710 140768
rect 1258 138336 218710 139200
rect 1258 136768 218710 137632
rect 1258 135225 218710 136064
rect 1258 135200 73213 135225
rect 1258 134471 68328 134496
rect 1258 133632 218710 134471
rect 1258 132903 137096 132928
rect 1258 132089 218710 132903
rect 1258 132064 65864 132089
rect 1258 131335 121416 131360
rect 1258 130521 218710 131335
rect 1258 130496 54552 130521
rect 1258 129767 61384 129792
rect 1258 128953 218710 129767
rect 1258 128928 46712 128953
rect 1258 128199 38269 128224
rect 1258 127385 218710 128199
rect 1258 127360 66895 127385
rect 1258 126631 44559 126656
rect 1258 125817 218710 126631
rect 1258 125792 45903 125817
rect 1258 125063 44396 125088
rect 1258 124249 218710 125063
rect 1258 124224 42117 124249
rect 1258 123495 40983 123520
rect 1258 122681 218710 123495
rect 1258 122656 39804 122681
rect 1258 121927 18221 121952
rect 1258 121113 218710 121927
rect 1258 121088 40588 121113
rect 1258 120359 11432 120384
rect 1258 119545 218710 120359
rect 1258 119520 24045 119545
rect 1258 118791 12733 118816
rect 1258 117977 218710 118791
rect 1258 117952 7245 117977
rect 1258 117223 41624 117248
rect 1258 116409 218710 117223
rect 1258 116384 6461 116409
rect 1258 115655 11949 115680
rect 1258 114841 218710 115655
rect 1258 114816 2989 114841
rect 1258 114087 18221 114112
rect 1258 113273 218710 114087
rect 1258 113248 14525 113273
rect 1258 112519 3437 112544
rect 1258 111705 218710 112519
rect 1258 111680 9037 111705
rect 1258 110951 58113 110976
rect 1258 110137 218710 110951
rect 1258 110112 15352 110137
rect 1258 109383 4445 109408
rect 1258 108569 218710 109383
rect 1258 108544 2989 108569
rect 1258 107815 3661 107840
rect 1258 107001 218710 107815
rect 1258 106976 47420 107001
rect 1258 106247 28568 106272
rect 1258 105433 218710 106247
rect 1258 105408 14301 105433
rect 1258 104679 3101 104704
rect 1258 103865 218710 104679
rect 1258 103840 7469 103865
rect 1258 103111 13517 103136
rect 1258 102297 218710 103111
rect 1258 102272 54427 102297
rect 1258 101543 20909 101568
rect 1258 100729 218710 101543
rect 1258 100704 18221 100729
rect 1258 99975 3101 100000
rect 1258 99161 218710 99975
rect 1258 99136 2989 99161
rect 1258 98407 6573 98432
rect 1258 97593 218710 98407
rect 1258 97568 50029 97593
rect 1258 96839 19453 96864
rect 1258 96025 218710 96839
rect 1258 96000 26173 96025
rect 1258 95271 68311 95296
rect 1258 94457 218710 95271
rect 1258 94432 45341 94457
rect 1258 93703 14142 93728
rect 1258 92889 218710 93703
rect 1258 92864 5798 92889
rect 1258 92135 4342 92160
rect 1258 91321 218710 92135
rect 1258 91296 14590 91321
rect 1258 90567 3567 90592
rect 1258 89753 218710 90567
rect 1258 89728 4118 89753
rect 1258 88999 15664 89024
rect 1258 88185 218710 88999
rect 1258 88160 30895 88185
rect 1258 87431 10390 87456
rect 1258 86617 218710 87431
rect 1258 86592 12462 86617
rect 1258 85863 55197 85888
rect 1258 85049 218710 85863
rect 1258 85024 9735 85049
rect 1258 84295 29766 84320
rect 1258 83481 218710 84295
rect 1258 83456 9847 83481
rect 1258 82727 27536 82752
rect 1258 81913 218710 82727
rect 1258 81888 5798 81913
rect 1258 81159 9718 81184
rect 1258 80345 218710 81159
rect 1258 80320 56231 80345
rect 1258 79591 3782 79616
rect 1258 78777 218710 79591
rect 1258 78752 31231 78777
rect 1258 78023 26014 78048
rect 1258 77209 218710 78023
rect 1258 77184 4006 77209
rect 1258 76455 36968 76480
rect 1258 75641 218710 76455
rect 1258 75616 9951 75641
rect 1258 74887 4566 74912
rect 1258 74073 218710 74887
rect 1258 74048 3903 74073
rect 1258 73319 36856 73344
rect 1258 72505 218710 73319
rect 1258 72480 24166 72505
rect 1258 71751 53096 71776
rect 1258 70937 218710 71751
rect 1258 70912 31032 70937
rect 1258 70183 51037 70208
rect 1258 69369 218710 70183
rect 1258 69344 15309 69369
rect 1258 68615 10381 68640
rect 1258 67801 218710 68615
rect 1258 67776 17437 67801
rect 1258 67047 10381 67072
rect 1258 66233 218710 67047
rect 1258 66208 10381 66233
rect 1258 65479 59885 65504
rect 1258 64665 218710 65479
rect 1258 64640 16205 64665
rect 1258 63911 45032 63936
rect 1258 63097 218710 63911
rect 1258 63072 17592 63097
rect 1258 62343 6461 62368
rect 1258 61529 218710 62343
rect 1258 61504 6461 61529
rect 1258 60775 59997 60800
rect 1258 59961 218710 60775
rect 1258 59936 23597 59961
rect 1258 59207 3885 59232
rect 1258 58393 218710 59207
rect 1258 58368 2989 58393
rect 1258 57639 11053 57664
rect 1258 56825 218710 57639
rect 1258 56800 31773 56825
rect 1258 56071 3997 56096
rect 1258 55257 218710 56071
rect 1258 55232 73549 55257
rect 1258 54503 33901 54528
rect 1258 53689 218710 54503
rect 1258 53664 18669 53689
rect 1258 52935 5789 52960
rect 1258 52121 218710 52935
rect 1258 52096 23933 52121
rect 1258 51367 6461 51392
rect 1258 50553 218710 51367
rect 1258 50528 6461 50553
rect 1258 49799 28413 49824
rect 1258 48985 218710 49799
rect 1258 48960 10829 48985
rect 1258 48231 6909 48256
rect 1258 47417 218710 48231
rect 1258 47392 73549 47417
rect 1258 46663 14637 46688
rect 1258 45849 218710 46663
rect 1258 45824 7917 45849
rect 1258 45095 20797 45120
rect 1258 44281 218710 45095
rect 1258 44256 10157 44281
rect 1258 43527 28637 43552
rect 1258 42713 218710 43527
rect 1258 42688 22141 42713
rect 1258 41959 14749 41984
rect 1258 41145 218710 41959
rect 1258 41120 22141 41145
rect 1258 40391 14232 40416
rect 1258 39577 218710 40391
rect 1258 39552 22701 39577
rect 1258 38823 29128 38848
rect 1258 38009 218710 38823
rect 1258 37984 29981 38009
rect 1258 37255 28861 37280
rect 1258 36441 218710 37255
rect 1258 36416 34349 36441
rect 1258 35687 34685 35712
rect 1258 34873 218710 35687
rect 1258 34848 56077 34873
rect 1258 34119 51149 34144
rect 1258 33305 218710 34119
rect 1258 33280 34125 33305
rect 1258 32551 34125 32576
rect 1258 31737 218710 32551
rect 1258 31712 41448 31737
rect 1258 30983 43912 31008
rect 1258 30169 218710 30983
rect 1258 30144 55336 30169
rect 1258 29415 83517 29440
rect 1258 28601 218710 29415
rect 1258 28576 63917 28601
rect 1258 27008 218710 27872
rect 1258 26279 74445 26304
rect 1258 25465 218710 26279
rect 1258 25440 62797 25465
rect 1258 23872 218710 24736
rect 1258 22329 218710 23168
rect 1258 22304 56792 22329
rect 1258 20736 218710 21600
rect 1258 19193 218710 20032
rect 1258 19168 89832 19193
rect 1258 18439 74109 18464
rect 1258 17600 218710 18439
rect 1258 16057 218710 16896
rect 1258 16032 93485 16057
rect 1258 14464 218710 15328
rect 1258 13735 77245 13760
rect 1258 12921 218710 13735
rect 1258 12896 49805 12921
rect 1258 11328 218710 12192
rect 1258 9760 218710 10624
rect 1258 8192 218710 9056
rect 1258 6624 218710 7488
rect 1258 5081 218710 5920
rect 1258 5056 32600 5081
rect 1258 4327 82397 4352
rect 1258 3488 218710 4327
<< pwell >>
rect 1258 156448 218710 156886
rect 1258 154880 218710 155584
rect 1258 153312 218710 154016
rect 1258 151744 218710 152448
rect 1258 150176 218710 150880
rect 1258 148608 218710 149312
rect 1258 147040 218710 147744
rect 1258 145472 218710 146176
rect 1258 143904 218710 144608
rect 1258 142336 218710 143040
rect 1258 140768 218710 141472
rect 1258 139200 218710 139904
rect 1258 137632 218710 138336
rect 1258 136064 218710 136768
rect 1258 134496 218710 135200
rect 1258 132928 218710 133632
rect 1258 131360 218710 132064
rect 1258 129792 218710 130496
rect 1258 128224 218710 128928
rect 1258 126656 218710 127360
rect 1258 125088 218710 125792
rect 1258 123520 218710 124224
rect 1258 121952 218710 122656
rect 1258 120384 218710 121088
rect 1258 118816 218710 119520
rect 1258 117248 218710 117952
rect 1258 115680 218710 116384
rect 1258 114112 218710 114816
rect 1258 112544 218710 113248
rect 1258 110976 218710 111680
rect 1258 109408 218710 110112
rect 1258 107840 218710 108544
rect 1258 106272 218710 106976
rect 1258 104704 218710 105408
rect 1258 103136 218710 103840
rect 1258 101568 218710 102272
rect 1258 100000 218710 100704
rect 1258 98432 218710 99136
rect 1258 96864 218710 97568
rect 1258 95296 218710 96000
rect 1258 93728 218710 94432
rect 1258 92160 218710 92864
rect 1258 90592 218710 91296
rect 1258 89024 218710 89728
rect 1258 87456 218710 88160
rect 1258 85888 218710 86592
rect 1258 84320 218710 85024
rect 1258 82752 218710 83456
rect 1258 81184 218710 81888
rect 1258 79616 218710 80320
rect 1258 78048 218710 78752
rect 1258 76480 218710 77184
rect 1258 74912 218710 75616
rect 1258 73344 218710 74048
rect 1258 71776 218710 72480
rect 1258 70208 218710 70912
rect 1258 68640 218710 69344
rect 1258 67072 218710 67776
rect 1258 65504 218710 66208
rect 1258 63936 218710 64640
rect 1258 62368 218710 63072
rect 1258 60800 218710 61504
rect 1258 59232 218710 59936
rect 1258 57664 218710 58368
rect 1258 56096 218710 56800
rect 1258 54528 218710 55232
rect 1258 52960 218710 53664
rect 1258 51392 218710 52096
rect 1258 49824 218710 50528
rect 1258 48256 218710 48960
rect 1258 46688 218710 47392
rect 1258 45120 218710 45824
rect 1258 43552 218710 44256
rect 1258 41984 218710 42688
rect 1258 40416 218710 41120
rect 1258 38848 218710 39552
rect 1258 37280 218710 37984
rect 1258 35712 218710 36416
rect 1258 34144 218710 34848
rect 1258 32576 218710 33280
rect 1258 31008 218710 31712
rect 1258 29440 218710 30144
rect 1258 27872 218710 28576
rect 1258 26304 218710 27008
rect 1258 24736 218710 25440
rect 1258 23168 218710 23872
rect 1258 21600 218710 22304
rect 1258 20032 218710 20736
rect 1258 18464 218710 19168
rect 1258 16896 218710 17600
rect 1258 15328 218710 16032
rect 1258 13760 218710 14464
rect 1258 12192 218710 12896
rect 1258 10624 218710 11328
rect 1258 9056 218710 9760
rect 1258 7488 218710 8192
rect 1258 5920 218710 6624
rect 1258 4352 218710 5056
rect 1258 3050 218710 3488
<< obsm1 >>
rect 1344 3076 218624 157218
<< metal2 >>
rect 8512 159200 8624 160000
rect 10304 159200 10416 160000
rect 12096 159200 12208 160000
rect 13888 159200 14000 160000
rect 15680 159200 15792 160000
rect 17472 159200 17584 160000
rect 19264 159200 19376 160000
rect 21056 159200 21168 160000
rect 22848 159200 22960 160000
rect 24640 159200 24752 160000
rect 26432 159200 26544 160000
rect 28224 159200 28336 160000
rect 30016 159200 30128 160000
rect 31808 159200 31920 160000
rect 33600 159200 33712 160000
rect 35392 159200 35504 160000
rect 37184 159200 37296 160000
rect 38976 159200 39088 160000
rect 40768 159200 40880 160000
rect 42560 159200 42672 160000
rect 44352 159200 44464 160000
rect 46144 159200 46256 160000
rect 47936 159200 48048 160000
rect 49728 159200 49840 160000
rect 51520 159200 51632 160000
rect 53312 159200 53424 160000
rect 55104 159200 55216 160000
rect 56896 159200 57008 160000
rect 58688 159200 58800 160000
rect 60480 159200 60592 160000
rect 62272 159200 62384 160000
rect 64064 159200 64176 160000
rect 65856 159200 65968 160000
rect 67648 159200 67760 160000
rect 69440 159200 69552 160000
rect 71232 159200 71344 160000
rect 73024 159200 73136 160000
rect 74816 159200 74928 160000
rect 76608 159200 76720 160000
rect 78400 159200 78512 160000
rect 80192 159200 80304 160000
rect 81984 159200 82096 160000
rect 83776 159200 83888 160000
rect 85568 159200 85680 160000
rect 87360 159200 87472 160000
rect 89152 159200 89264 160000
rect 90944 159200 91056 160000
rect 92736 159200 92848 160000
rect 94528 159200 94640 160000
rect 96320 159200 96432 160000
rect 98112 159200 98224 160000
rect 99904 159200 100016 160000
rect 101696 159200 101808 160000
rect 103488 159200 103600 160000
rect 105280 159200 105392 160000
rect 107072 159200 107184 160000
rect 108864 159200 108976 160000
rect 110656 159200 110768 160000
rect 112448 159200 112560 160000
rect 114240 159200 114352 160000
rect 116032 159200 116144 160000
rect 117824 159200 117936 160000
rect 119616 159200 119728 160000
rect 121408 159200 121520 160000
rect 123200 159200 123312 160000
rect 124992 159200 125104 160000
rect 126784 159200 126896 160000
rect 128576 159200 128688 160000
rect 130368 159200 130480 160000
rect 132160 159200 132272 160000
rect 133952 159200 134064 160000
rect 135744 159200 135856 160000
rect 137536 159200 137648 160000
rect 139328 159200 139440 160000
rect 141120 159200 141232 160000
rect 142912 159200 143024 160000
rect 144704 159200 144816 160000
rect 146496 159200 146608 160000
rect 148288 159200 148400 160000
rect 150080 159200 150192 160000
rect 151872 159200 151984 160000
rect 153664 159200 153776 160000
rect 155456 159200 155568 160000
rect 157248 159200 157360 160000
rect 159040 159200 159152 160000
rect 160832 159200 160944 160000
rect 162624 159200 162736 160000
rect 164416 159200 164528 160000
rect 166208 159200 166320 160000
rect 168000 159200 168112 160000
rect 169792 159200 169904 160000
rect 171584 159200 171696 160000
rect 173376 159200 173488 160000
rect 175168 159200 175280 160000
rect 176960 159200 177072 160000
rect 178752 159200 178864 160000
rect 180544 159200 180656 160000
rect 182336 159200 182448 160000
rect 184128 159200 184240 160000
rect 185920 159200 186032 160000
rect 187712 159200 187824 160000
rect 189504 159200 189616 160000
rect 191296 159200 191408 160000
rect 193088 159200 193200 160000
rect 194880 159200 194992 160000
rect 196672 159200 196784 160000
rect 198464 159200 198576 160000
rect 200256 159200 200368 160000
rect 202048 159200 202160 160000
rect 203840 159200 203952 160000
rect 205632 159200 205744 160000
rect 207424 159200 207536 160000
rect 209216 159200 209328 160000
rect 211008 159200 211120 160000
rect 2240 0 2352 800
rect 5600 0 5712 800
rect 8960 0 9072 800
rect 12320 0 12432 800
rect 15680 0 15792 800
rect 19040 0 19152 800
rect 22400 0 22512 800
rect 25760 0 25872 800
rect 29120 0 29232 800
rect 32480 0 32592 800
rect 35840 0 35952 800
rect 39200 0 39312 800
rect 42560 0 42672 800
rect 45920 0 46032 800
rect 49280 0 49392 800
rect 52640 0 52752 800
rect 56000 0 56112 800
rect 59360 0 59472 800
rect 62720 0 62832 800
rect 66080 0 66192 800
rect 69440 0 69552 800
rect 72800 0 72912 800
rect 76160 0 76272 800
rect 79520 0 79632 800
rect 82880 0 82992 800
rect 86240 0 86352 800
rect 89600 0 89712 800
rect 92960 0 93072 800
rect 96320 0 96432 800
rect 99680 0 99792 800
rect 103040 0 103152 800
rect 106400 0 106512 800
rect 109760 0 109872 800
rect 113120 0 113232 800
rect 116480 0 116592 800
rect 119840 0 119952 800
rect 123200 0 123312 800
rect 126560 0 126672 800
rect 129920 0 130032 800
rect 133280 0 133392 800
rect 136640 0 136752 800
rect 140000 0 140112 800
rect 143360 0 143472 800
rect 146720 0 146832 800
rect 150080 0 150192 800
rect 153440 0 153552 800
rect 156800 0 156912 800
rect 160160 0 160272 800
rect 163520 0 163632 800
rect 166880 0 166992 800
rect 170240 0 170352 800
rect 173600 0 173712 800
rect 176960 0 177072 800
rect 180320 0 180432 800
rect 183680 0 183792 800
rect 187040 0 187152 800
rect 190400 0 190512 800
rect 193760 0 193872 800
rect 197120 0 197232 800
rect 200480 0 200592 800
rect 203840 0 203952 800
rect 207200 0 207312 800
rect 210560 0 210672 800
rect 213920 0 214032 800
rect 217280 0 217392 800
<< obsm2 >>
rect 1596 159140 8452 159348
rect 8684 159140 10244 159348
rect 10476 159140 12036 159348
rect 12268 159140 13828 159348
rect 14060 159140 15620 159348
rect 15852 159140 17412 159348
rect 17644 159140 19204 159348
rect 19436 159140 20996 159348
rect 21228 159140 22788 159348
rect 23020 159140 24580 159348
rect 24812 159140 26372 159348
rect 26604 159140 28164 159348
rect 28396 159140 29956 159348
rect 30188 159140 31748 159348
rect 31980 159140 33540 159348
rect 33772 159140 35332 159348
rect 35564 159140 37124 159348
rect 37356 159140 38916 159348
rect 39148 159140 40708 159348
rect 40940 159140 42500 159348
rect 42732 159140 44292 159348
rect 44524 159140 46084 159348
rect 46316 159140 47876 159348
rect 48108 159140 49668 159348
rect 49900 159140 51460 159348
rect 51692 159140 53252 159348
rect 53484 159140 55044 159348
rect 55276 159140 56836 159348
rect 57068 159140 58628 159348
rect 58860 159140 60420 159348
rect 60652 159140 62212 159348
rect 62444 159140 64004 159348
rect 64236 159140 65796 159348
rect 66028 159140 67588 159348
rect 67820 159140 69380 159348
rect 69612 159140 71172 159348
rect 71404 159140 72964 159348
rect 73196 159140 74756 159348
rect 74988 159140 76548 159348
rect 76780 159140 78340 159348
rect 78572 159140 80132 159348
rect 80364 159140 81924 159348
rect 82156 159140 83716 159348
rect 83948 159140 85508 159348
rect 85740 159140 87300 159348
rect 87532 159140 89092 159348
rect 89324 159140 90884 159348
rect 91116 159140 92676 159348
rect 92908 159140 94468 159348
rect 94700 159140 96260 159348
rect 96492 159140 98052 159348
rect 98284 159140 99844 159348
rect 100076 159140 101636 159348
rect 101868 159140 103428 159348
rect 103660 159140 105220 159348
rect 105452 159140 107012 159348
rect 107244 159140 108804 159348
rect 109036 159140 110596 159348
rect 110828 159140 112388 159348
rect 112620 159140 114180 159348
rect 114412 159140 115972 159348
rect 116204 159140 117764 159348
rect 117996 159140 119556 159348
rect 119788 159140 121348 159348
rect 121580 159140 123140 159348
rect 123372 159140 124932 159348
rect 125164 159140 126724 159348
rect 126956 159140 128516 159348
rect 128748 159140 130308 159348
rect 130540 159140 132100 159348
rect 132332 159140 133892 159348
rect 134124 159140 135684 159348
rect 135916 159140 137476 159348
rect 137708 159140 139268 159348
rect 139500 159140 141060 159348
rect 141292 159140 142852 159348
rect 143084 159140 144644 159348
rect 144876 159140 146436 159348
rect 146668 159140 148228 159348
rect 148460 159140 150020 159348
rect 150252 159140 151812 159348
rect 152044 159140 153604 159348
rect 153836 159140 155396 159348
rect 155628 159140 157188 159348
rect 157420 159140 158980 159348
rect 159212 159140 160772 159348
rect 161004 159140 162564 159348
rect 162796 159140 164356 159348
rect 164588 159140 166148 159348
rect 166380 159140 167940 159348
rect 168172 159140 169732 159348
rect 169964 159140 171524 159348
rect 171756 159140 173316 159348
rect 173548 159140 175108 159348
rect 175340 159140 176900 159348
rect 177132 159140 178692 159348
rect 178924 159140 180484 159348
rect 180716 159140 182276 159348
rect 182508 159140 184068 159348
rect 184300 159140 185860 159348
rect 186092 159140 187652 159348
rect 187884 159140 189444 159348
rect 189676 159140 191236 159348
rect 191468 159140 193028 159348
rect 193260 159140 194820 159348
rect 195052 159140 196612 159348
rect 196844 159140 198404 159348
rect 198636 159140 200196 159348
rect 200428 159140 201988 159348
rect 202220 159140 203780 159348
rect 204012 159140 205572 159348
rect 205804 159140 207364 159348
rect 207596 159140 209156 159348
rect 209388 159140 210948 159348
rect 211180 159140 217588 159348
rect 1596 860 217588 159140
rect 1596 700 2180 860
rect 2412 700 5540 860
rect 5772 700 8900 860
rect 9132 700 12260 860
rect 12492 700 15620 860
rect 15852 700 18980 860
rect 19212 700 22340 860
rect 22572 700 25700 860
rect 25932 700 29060 860
rect 29292 700 32420 860
rect 32652 700 35780 860
rect 36012 700 39140 860
rect 39372 700 42500 860
rect 42732 700 45860 860
rect 46092 700 49220 860
rect 49452 700 52580 860
rect 52812 700 55940 860
rect 56172 700 59300 860
rect 59532 700 62660 860
rect 62892 700 66020 860
rect 66252 700 69380 860
rect 69612 700 72740 860
rect 72972 700 76100 860
rect 76332 700 79460 860
rect 79692 700 82820 860
rect 83052 700 86180 860
rect 86412 700 89540 860
rect 89772 700 92900 860
rect 93132 700 96260 860
rect 96492 700 99620 860
rect 99852 700 102980 860
rect 103212 700 106340 860
rect 106572 700 109700 860
rect 109932 700 113060 860
rect 113292 700 116420 860
rect 116652 700 119780 860
rect 120012 700 123140 860
rect 123372 700 126500 860
rect 126732 700 129860 860
rect 130092 700 133220 860
rect 133452 700 136580 860
rect 136812 700 139940 860
rect 140172 700 143300 860
rect 143532 700 146660 860
rect 146892 700 150020 860
rect 150252 700 153380 860
rect 153612 700 156740 860
rect 156972 700 160100 860
rect 160332 700 163460 860
rect 163692 700 166820 860
rect 167052 700 170180 860
rect 170412 700 173540 860
rect 173772 700 176900 860
rect 177132 700 180260 860
rect 180492 700 183620 860
rect 183852 700 186980 860
rect 187212 700 190340 860
rect 190572 700 193700 860
rect 193932 700 197060 860
rect 197292 700 200420 860
rect 200652 700 203780 860
rect 204012 700 207140 860
rect 207372 700 210500 860
rect 210732 700 213860 860
rect 214092 700 217220 860
rect 217452 700 217588 860
<< obsm3 >>
rect 1586 3108 204430 158452
<< metal4 >>
rect 4448 3076 4768 156860
rect 19808 3076 20128 156860
rect 35168 3076 35488 156860
rect 50528 3076 50848 156860
rect 65888 3076 66208 156860
rect 81248 3076 81568 156860
rect 96608 3076 96928 156860
rect 111968 3076 112288 156860
rect 127328 3076 127648 156860
rect 142688 3076 143008 156860
rect 158048 3076 158368 156860
rect 173408 3076 173728 156860
rect 188768 3076 189088 156860
rect 204128 3076 204448 156860
<< obsm4 >>
rect 7084 156920 166404 158350
rect 7084 11106 19748 156920
rect 20188 11106 35108 156920
rect 35548 11106 50468 156920
rect 50908 11106 65828 156920
rect 66268 11106 81188 156920
rect 81628 11106 96548 156920
rect 96988 11106 111908 156920
rect 112348 11106 127268 156920
rect 127708 11106 142628 156920
rect 143068 11106 157988 156920
rect 158428 11106 166404 156920
<< labels >>
rlabel metal2 s 8512 159200 8624 160000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 62272 159200 62384 160000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 67648 159200 67760 160000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 73024 159200 73136 160000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 78400 159200 78512 160000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 83776 159200 83888 160000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 89152 159200 89264 160000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 94528 159200 94640 160000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 99904 159200 100016 160000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 105280 159200 105392 160000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 110656 159200 110768 160000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 13888 159200 14000 160000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 116032 159200 116144 160000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 121408 159200 121520 160000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 126784 159200 126896 160000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 132160 159200 132272 160000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 137536 159200 137648 160000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 142912 159200 143024 160000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 148288 159200 148400 160000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 153664 159200 153776 160000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 159040 159200 159152 160000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 164416 159200 164528 160000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 19264 159200 19376 160000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 169792 159200 169904 160000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 175168 159200 175280 160000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 180544 159200 180656 160000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 185920 159200 186032 160000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 191296 159200 191408 160000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 196672 159200 196784 160000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 202048 159200 202160 160000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 207424 159200 207536 160000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 24640 159200 24752 160000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 30016 159200 30128 160000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35392 159200 35504 160000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 40768 159200 40880 160000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 46144 159200 46256 160000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 51520 159200 51632 160000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 56896 159200 57008 160000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 10304 159200 10416 160000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 64064 159200 64176 160000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 69440 159200 69552 160000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 74816 159200 74928 160000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 80192 159200 80304 160000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 85568 159200 85680 160000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 90944 159200 91056 160000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 96320 159200 96432 160000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 101696 159200 101808 160000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 107072 159200 107184 160000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 112448 159200 112560 160000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15680 159200 15792 160000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 117824 159200 117936 160000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 123200 159200 123312 160000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 128576 159200 128688 160000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 133952 159200 134064 160000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 139328 159200 139440 160000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 144704 159200 144816 160000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 150080 159200 150192 160000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 155456 159200 155568 160000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 160832 159200 160944 160000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 166208 159200 166320 160000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 21056 159200 21168 160000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 171584 159200 171696 160000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 176960 159200 177072 160000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 182336 159200 182448 160000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 187712 159200 187824 160000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 193088 159200 193200 160000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 198464 159200 198576 160000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 203840 159200 203952 160000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 209216 159200 209328 160000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26432 159200 26544 160000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 31808 159200 31920 160000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 37184 159200 37296 160000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 42560 159200 42672 160000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 47936 159200 48048 160000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 53312 159200 53424 160000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 58688 159200 58800 160000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 12096 159200 12208 160000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 65856 159200 65968 160000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 71232 159200 71344 160000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 76608 159200 76720 160000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 81984 159200 82096 160000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 87360 159200 87472 160000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 92736 159200 92848 160000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 98112 159200 98224 160000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 103488 159200 103600 160000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 108864 159200 108976 160000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 114240 159200 114352 160000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 17472 159200 17584 160000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 119616 159200 119728 160000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 124992 159200 125104 160000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 130368 159200 130480 160000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 135744 159200 135856 160000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 141120 159200 141232 160000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 146496 159200 146608 160000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 151872 159200 151984 160000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 157248 159200 157360 160000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 162624 159200 162736 160000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 168000 159200 168112 160000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 22848 159200 22960 160000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 173376 159200 173488 160000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 178752 159200 178864 160000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 184128 159200 184240 160000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 189504 159200 189616 160000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 194880 159200 194992 160000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 200256 159200 200368 160000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 205632 159200 205744 160000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 211008 159200 211120 160000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 28224 159200 28336 160000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 33600 159200 33712 160000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 38976 159200 39088 160000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 44352 159200 44464 160000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 49728 159200 49840 160000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 55104 159200 55216 160000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 60480 159200 60592 160000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 5600 0 5712 800 6 la_data_out[0]
port 115 nsew signal output
rlabel metal2 s 39200 0 39312 800 6 la_data_out[10]
port 116 nsew signal output
rlabel metal2 s 42560 0 42672 800 6 la_data_out[11]
port 117 nsew signal output
rlabel metal2 s 45920 0 46032 800 6 la_data_out[12]
port 118 nsew signal output
rlabel metal2 s 49280 0 49392 800 6 la_data_out[13]
port 119 nsew signal output
rlabel metal2 s 52640 0 52752 800 6 la_data_out[14]
port 120 nsew signal output
rlabel metal2 s 56000 0 56112 800 6 la_data_out[15]
port 121 nsew signal output
rlabel metal2 s 59360 0 59472 800 6 la_data_out[16]
port 122 nsew signal output
rlabel metal2 s 62720 0 62832 800 6 la_data_out[17]
port 123 nsew signal output
rlabel metal2 s 66080 0 66192 800 6 la_data_out[18]
port 124 nsew signal output
rlabel metal2 s 69440 0 69552 800 6 la_data_out[19]
port 125 nsew signal output
rlabel metal2 s 8960 0 9072 800 6 la_data_out[1]
port 126 nsew signal output
rlabel metal2 s 72800 0 72912 800 6 la_data_out[20]
port 127 nsew signal output
rlabel metal2 s 76160 0 76272 800 6 la_data_out[21]
port 128 nsew signal output
rlabel metal2 s 79520 0 79632 800 6 la_data_out[22]
port 129 nsew signal output
rlabel metal2 s 82880 0 82992 800 6 la_data_out[23]
port 130 nsew signal output
rlabel metal2 s 86240 0 86352 800 6 la_data_out[24]
port 131 nsew signal output
rlabel metal2 s 89600 0 89712 800 6 la_data_out[25]
port 132 nsew signal output
rlabel metal2 s 92960 0 93072 800 6 la_data_out[26]
port 133 nsew signal output
rlabel metal2 s 96320 0 96432 800 6 la_data_out[27]
port 134 nsew signal output
rlabel metal2 s 99680 0 99792 800 6 la_data_out[28]
port 135 nsew signal output
rlabel metal2 s 103040 0 103152 800 6 la_data_out[29]
port 136 nsew signal output
rlabel metal2 s 12320 0 12432 800 6 la_data_out[2]
port 137 nsew signal output
rlabel metal2 s 106400 0 106512 800 6 la_data_out[30]
port 138 nsew signal output
rlabel metal2 s 109760 0 109872 800 6 la_data_out[31]
port 139 nsew signal output
rlabel metal2 s 113120 0 113232 800 6 la_data_out[32]
port 140 nsew signal output
rlabel metal2 s 116480 0 116592 800 6 la_data_out[33]
port 141 nsew signal output
rlabel metal2 s 119840 0 119952 800 6 la_data_out[34]
port 142 nsew signal output
rlabel metal2 s 123200 0 123312 800 6 la_data_out[35]
port 143 nsew signal output
rlabel metal2 s 126560 0 126672 800 6 la_data_out[36]
port 144 nsew signal output
rlabel metal2 s 129920 0 130032 800 6 la_data_out[37]
port 145 nsew signal output
rlabel metal2 s 133280 0 133392 800 6 la_data_out[38]
port 146 nsew signal output
rlabel metal2 s 136640 0 136752 800 6 la_data_out[39]
port 147 nsew signal output
rlabel metal2 s 15680 0 15792 800 6 la_data_out[3]
port 148 nsew signal output
rlabel metal2 s 140000 0 140112 800 6 la_data_out[40]
port 149 nsew signal output
rlabel metal2 s 143360 0 143472 800 6 la_data_out[41]
port 150 nsew signal output
rlabel metal2 s 146720 0 146832 800 6 la_data_out[42]
port 151 nsew signal output
rlabel metal2 s 150080 0 150192 800 6 la_data_out[43]
port 152 nsew signal output
rlabel metal2 s 153440 0 153552 800 6 la_data_out[44]
port 153 nsew signal output
rlabel metal2 s 156800 0 156912 800 6 la_data_out[45]
port 154 nsew signal output
rlabel metal2 s 160160 0 160272 800 6 la_data_out[46]
port 155 nsew signal output
rlabel metal2 s 163520 0 163632 800 6 la_data_out[47]
port 156 nsew signal output
rlabel metal2 s 166880 0 166992 800 6 la_data_out[48]
port 157 nsew signal output
rlabel metal2 s 170240 0 170352 800 6 la_data_out[49]
port 158 nsew signal output
rlabel metal2 s 19040 0 19152 800 6 la_data_out[4]
port 159 nsew signal output
rlabel metal2 s 173600 0 173712 800 6 la_data_out[50]
port 160 nsew signal output
rlabel metal2 s 176960 0 177072 800 6 la_data_out[51]
port 161 nsew signal output
rlabel metal2 s 180320 0 180432 800 6 la_data_out[52]
port 162 nsew signal output
rlabel metal2 s 183680 0 183792 800 6 la_data_out[53]
port 163 nsew signal output
rlabel metal2 s 187040 0 187152 800 6 la_data_out[54]
port 164 nsew signal output
rlabel metal2 s 190400 0 190512 800 6 la_data_out[55]
port 165 nsew signal output
rlabel metal2 s 193760 0 193872 800 6 la_data_out[56]
port 166 nsew signal output
rlabel metal2 s 197120 0 197232 800 6 la_data_out[57]
port 167 nsew signal output
rlabel metal2 s 200480 0 200592 800 6 la_data_out[58]
port 168 nsew signal output
rlabel metal2 s 203840 0 203952 800 6 la_data_out[59]
port 169 nsew signal output
rlabel metal2 s 22400 0 22512 800 6 la_data_out[5]
port 170 nsew signal output
rlabel metal2 s 207200 0 207312 800 6 la_data_out[60]
port 171 nsew signal output
rlabel metal2 s 210560 0 210672 800 6 la_data_out[61]
port 172 nsew signal output
rlabel metal2 s 213920 0 214032 800 6 la_data_out[62]
port 173 nsew signal output
rlabel metal2 s 217280 0 217392 800 6 la_data_out[63]
port 174 nsew signal output
rlabel metal2 s 25760 0 25872 800 6 la_data_out[6]
port 175 nsew signal output
rlabel metal2 s 29120 0 29232 800 6 la_data_out[7]
port 176 nsew signal output
rlabel metal2 s 32480 0 32592 800 6 la_data_out[8]
port 177 nsew signal output
rlabel metal2 s 35840 0 35952 800 6 la_data_out[9]
port 178 nsew signal output
rlabel metal4 s 4448 3076 4768 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 156860 6 vdd
port 179 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 156860 6 vss
port 180 nsew ground bidirectional
rlabel metal2 s 2240 0 2352 800 6 wb_clk_i
port 181 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 220000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16001752
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/wrapped_as2650/runs/23_11_01_11_20/results/signoff/wrapped_as2650.magic.gds
string GDS_START 536280
<< end >>

